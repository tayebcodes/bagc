PK   ���X�8lѷ  �-    cirkitFile.json�]�nc7�~���f��K�Kz2� I�'���H7�[Z;n�+��d�<о�>��d�\t�������D>�,Y�UE��o�e����(����jy3_\M^r=�|��Sh?e�����b���i�?L^���V�^WY��x����V�E��Ϥ�]��Zg��2����r#/�����.h�%���Ug��V�Ъ[ZuG��i�9q�9���[N.'"��ǉ��D���]��jS�<���F����ȸѹ.��3�Y����D�
��%BW�+Ԙ��ބ:�W �Rf�y�9W�E-+� ���e�xeBpY����FAݐgU���̎խ�7eaEf���]�g9�nP*��{��X]Q�<��C?����|BVU��L�Zu)å)�EB�0#M�zMkڎ4�'�����Z��I'j��k����
ʱ�׬t��؂�Oш��%Q�I�F�T#���$q1���XcI\��[�[G�:r9!4�IM[J�b��J1��Y.����J�����*�ƨr|�bZ���G�#�履��ל�Y�57�u�J�:7�Υe%i-������F�����%�Ҵ�4=�nQ�J�Ng%�P9@���8�`@E�h�=�nT�cC�|t�Z>	����)Ѝ�m)MkJ�c�fFV!x���r�x����C�s�R�6�c�F�<�1T�'A7��Ӡ�1��8?��	��1tk��R��ɠB�xM��B4�A)UyE�1t�Z���1tKŌS�τP P�3E�PeT�qk���Q-��95�M���E.u��M*����yw����1nRZkܤ��2RZ��I}�#-#BB�l��H����X��n!<9�g��@hy��H㑠����4	-�����B~��EEdGM
�.�m���9\$�2b��Ga�C��=�P,.K�ф�g��7��"O($�"�PQI��$Tt*&	���KB�'������<�$�ifO3x�4�i0��s42iP,ҠX$��iP,ҠX4(�k/mE!�Fq��0���돝�`�S�4(��1(d�ؑ�!nP����k�ڝ�2�e"�$�e],��b�F�4�X6(����r����DnZO>�u(���\�R\��µ�D��y^�"'�: #�~�~��z�|f�,%�Gr�#&|I�{�v{s���[��e��uܿ�b7#/VI����*G�rPF�M�2Bn��r�l���n��q	��FF�p�1A��S�[�#{'ح&��	3�w��F�%�ُ݊:����q�nU���~�`������Ɔ�����0���r߿a����.6~@�"����l�y���������m���7����qܫ�v���8.��LBE%�P�I��$Tl*.	��
O#$�f�4����<�4�i��@���0Ob��"�E"M��"�E�4(iP,ҠX�A�H�b��2�e"�$�e�4(�iP,ӠXF16�K�r|�8.��a�a�t*����ҩ�:�K�rPF�8.��A��t*e���ҩ�:�K�rXF�8.��aa�t*�e���ҩ�:�K�rPF�8.��A^�q\:�����t*��ǥS9�:�K�rX�`�t*yA�q�Tڼ�>����֧q/��/��BO'�������2Uy1��X,�j9y���c�Ѿ�&3�A�̙�Yb)��k���Kځ>R��e��y���5�eJ>q���W����4��Zƍ�	Z�\Z#�6nN� �g��8�26�G�HHMRP�M��D�.:?Z�)ꄝ�id�M����5:��	d��G�F�W'X:���c)p�M�'�\RF��hQZF��O�m��)-�䌌 Q�$��i'�FZFFT(�;J�G�Pt>��vJ���򈳁�+���Gg�J�`���Q��S�X��i'Ǵ'.>D�s��k#F�t�x���X����4�����ZF��"�;��IM�ç���ĦGp��5�OL���L�O:�x�����n�aY}\�\��ܵ�#����?ږ���:�'c �3@ܧ8XO�d`@�F�D�ݚs�|L���;ED�=���3��R�;g�ow������3+��d��|�Pq�,��l�&���_;.�'r�_H#��q���	8 �XN���?� ���v���x@���rp�g:č��c��d$q:ϱ}2���D��a��cs�iX���$��{�t�[�{8��=}�����3��� n��@�aW�� qs����������3����sl�Ӈ���O4I�i�Op��������g	_|F7MRy�'>҆!�r��43����A���4I"@�#8�����8⁜q�g��ĳXI�H<����%�F�N�Y��B8�Q��Y��Q�g�²��_mSqn�^ܥ�y:o�%5K�e��Kb}E�ψ�5��!ַ���X��s� 8��
aN�0���SQȩ0�T6�3Y��kG��$)6*0Y�R�)��l�dv��F�Z�l�=z$��鑎H�!��(">�f����茚=z#�&>�&i��b\��*�%U�J��T�+��W��I2�z�-9�i3{���I)��hg���~�G���v�d�96{�(;�;$K�n�dGw���7q�E���I��'Ytf�9Jdr�d)�;vH�2vxɢ�w"%�M㉔,6�g���a`lb����`3|�ȍſ��>{�F�t�����tP���@qc���;t�P�ЙBq�C��R�QйC{�F��!�����Η`�YtZ�����ȍicl��9���vp72�ЩG{��6頳�O'�d�e�Z���Ƹ'��?N�\������`�B�]����ӯAy3sD5(m�Ј����x�ќ��XC��NZs٤���/o�u��k�XC6,�2֐���5d�!��	�h�=l��2^ٚ`lý0&�^9/KD�ٲ�A�PԶP���*��N� �d)4LhJ�J��<4��_�6���ؔ��ZC�2���/2W� �ш��VڭKb�ٽ�c��{�0�N�
��S��;0j�S��:0ʧS�:rW��T�U�����r��,f�R\�P|9���H �L)@�/��sE�'�� ����6&�P��,�}�x^C��������"�"3U�*9��e���)�`h�o��,�4�HX�kV����KTm�%W�ec	=r0�����HS°u�.��c��:��4�&�U�1[�V�z31jSiⲾ�A#�����JՁi��f�D� �u� }�L�`Z�P�D_Z Rmz�j���nW���K���d���2/Mь'(�۵~��VQ=_��޿(VB��d��$n�IP���7'��Gͳ9tw����(�H�n���`����2�'$]������.CQ�t�A0��D�=9t�	�P�Q]��̜%C�Ё'�5i��_'�$�<��X�jj�a���W��.�q3��ðA�Rsb�&f�i2�A��H�77����ɏ���(��=]��qL��_Yŏ�\����nKO��׷��E���yŇ������Wr�Jm^��+�y��������Wv��m^��+�y����h��p��pǃߍ�>~7"|8$�nH�pL�]�������|�u~7���.//�%���",c��zqq9�Ym�o�h��KXE����ћ��Z��U�^����|5_\A��L0�8�*�g��f
(EpUS�V��[�1�J�ݗU�t^�`X^���-�P-o�b:�_ݬ�U�!�	�N'����5{���H{�,.�M�~4���T+�~z�[��߼����6k�ؾQ��5����U�h=��ϥ�.]�i=׭��\��������Z��yތC�Kn���3v�l����>��gj�Ll��g�5�����>��gr�Ll���g�&6{�������m9_lq3�39�0bWp?s�;��o�IhXͬҙ6�K4�\	���3%��r˫L3���*�l'�yØ�8ò��x��&�����%���͌o��0�z�ȍ+>��N�;3��;�gJu�I���1ߩ���SHgjN+ԎZ8F�΄���2=Q�ݒҍ��Sv��t#�>���L#�!��(c�.��Hr�j��#�R��oV���O0XW�c����t�s���O~������͋>���/�����O�ײ��������U��˰��~m��>�6�z�i!�p�To>,>��6�'/�pyS��N�����;ܼ����>�ٶ�Tn���O���U�*~w���=3�2����n����}��ס��|W#w�����9�����kt��^\����U�}�%*�Aj��Z��Z��]���������Sf� s�K.�T�V��Rf��`ⴕ��N�}��g%��ы�uJZw60J��xX�m�����7_��>O��i��������E�z��~̬��p���ܞd������4��W_?���Y�X�,R+�u\���lb��o.֟f�b�לf��|a�L�n��m���W�	��;/s�y�3^� ދ�Y��ȡ�gU��c��s`�p�v-Y�����q��|�9�r�g��J��]G��S�b���k7㦂�;OT���ޙ��6���tSe7ަ�4s�u�-7�Z!�����[B���m1�
�b#� x��$�X
t�d Ä�f���f���fڂ1�z�iW�Li�`�s�q�]�[�+eP�A����	LM���-?5�7e���Цs�lZ�ܨYtcTK`-5�( P�t�Y�o�"U�8c��y�5�)BL�4Gg���N���FM9��=,��8i$̒Mkq��`�ʻ�x{��CϹ��(]��e��N�0����:W���i���n�	�KY�!=`��	��X!ܝ�VS	��j�����$3y&�ہR\�Y�W�D
PѹB�#�)b31�u|z������';	Y�t�P'n6f�݂]/�X2I�lcf��c��l�Pǎ6jڏ M�.���`L0$��SX���ߙ	�Fh�b�m c��U�LSy�C�jo��-���Ԉ��"nw�w����ct�]~�@����~����_���۷��{�����sz��)ɬ��	���T��N��g��Mu��t�l�=�EȾ�n�kVZ�Z.n���~l[�Zr����Oo&�'N"A�y�]��)�B6/�r��m��"xO�|����}n��r��ꞟ�R���CtG禹E�o|�f|���淈�Y����(T�ٷ�s�����᪼��_�l���j���~��W���hEa���8.�Sxq:h��d�8d��`�ZfY��)��9���5����~�,�����npa�e�[mTǾ����,˲�:J+]�Ns��-Pw��!��i�3]���T���uNXfA���zP\���ycA��g��7�)A�C���
����/���:�<�<sB>�9�� ��C�)75R�LB��k�4NbO�n�CS5g��Nr�A�Z�-��1PS�Ie\�7bu(U�UV�����xp�gK��>ap��0���RT_|��o���z�����?�ʮ����g����Ϊ���`3�`��+��S���G?&�V`��Dm�.\?�Ig��
F���o~���y�>O��Z�ͬ��9Iǧ�����x.��4QTփ'4]�y���_~�<;�x��1C�B����{���O��3c�Bj�cޞ�p,*+���|���٩f�ig��JI�LsvIi�$,m�Z}�ى���<;�g���l�N/�{l<�3��!�4�-*�}z��<c��� �O�Lx0ځ�eU�1ʸW3�A#��O�r�!�7�̬X'�P���r-��h����K��-�0�E(>T����o��j�����?@��o�`� a�&/��*0"����苰��w�Uټzpn��XuU�%����Z�OoS���L���b+�>4�~{���$�]��/�6Z�&>}�c���(��)�����X`ڔ��D����u�m[Jw.^�(���w��L=h0]K��.QZBh<4��-4Lh4��w�t��,�1����e@B��.!4,G�64�n}�X����R(�1(� �����#x{lh��\p-v��'t\��Ј�^�Jik(4p��
��#�;������w�f��m��R�#q\���ƠP���J�\b�G���=%�t/7�a���x�B���#�����ʕ���qX<�"�;vA: %�����n��!��@��3�<嚥���x��I�{��Q|�[��$��
�w�cT!���
%@���D�49eI4��b&Q���-$w#��a����~]qkOIW�oV�8�PR]��-s�D.�7
���xT�Gpw$*�q/�v����aT)��r�&k��j�9F�	N�"%zp�+.	|b��m�#�;=�v�E��=.Dc�R���X'���GvJ��P�
�\��t�x��Z*􈇠Gu��<�f����d|��ny��N)��B&�wZm!��i"v�H�)p���@�Ȇ�=vu�}�!�r���`-�� yǬm���m�f�A2c�H[�J톅n.ܤ�EB���k�`� �߃�;uz�}@fg����]��<y<ǘ/Sz�ܗW{��#�{�ۚ��c��P�EfP��a�G��R&n�t�H�Ia��Fw�6��v��R|�&�JUh�y�>x��E�ڪ ���}hg���w���a�R<w�I��#�gb�R���*�H������;,x��0�WH�EwqC�B��u�%:����(���}E4����=���Bk����8��ǗR�C���F�R)�����#A�ۓ��HD�'t\�G��cÏ�#x{RА(}�+����}�q�qoO
��Y�"ʐ��}�3�8^�G�L��!�����8�P�%�������,L��&�}�5!0����d�������s�\_j$�чƠ�ӂ�û���#�;	0⩝�Ku�C(5��9�b���q:���XL��-���ZL��h�0���3�@�54������������py3y�r��1�WU~�n����_���7�C�#��������_��b9��\0���PK   ���X��2i  �t  /   images/0d24f7ca-0a17-4a90-9ee7-368ce6dafe9a.png�uTTm�>< HI�tw-�t9tJ�tw�����JK�  �-����x��}����[���[�c�^{��W�u��y�ᕺ�<&:):�TT���a ��C�N�s��^n'-��(-M���lm��
Rx�����4��{[�2�mHHru&HSJ
M֯�('�\�Hׅ�0��k��0K�(Z""�|=bK��a��MTO�gW��g�~}1]��=��vc�."Od&y�B-�F�u�V +';�BBK�>����4Gzx� �2�����R�����<�eE&1���"�EŻ�.<�kG{{FڦW�@�i�l�m|��[�<���Gô�-Ee��G-"P��x0
R��6�yN���J7���ĊmF��
�AU�(�aP��3oW�p{���%��[?�C����6���P����#�����EjJ�)�`/���>�7����2,��y��}��Vx8h�
���T����R;E}g�j��O�}Zg�E��x=�^�wU��;���(N�G�P�T�j`�f�{Y6ב[v�&���҅i/�3�Sk�p?��w�\��: 	ɣ�U�+���7����85�>ggo1��D*�ZS�98�`t@\}�)eOZ��ai�X�(5���^l��,��G�Y�#��<�qK�\���z �LU���-�K����0��é�w>�?Z�\�(}W�N��I'6p#�K���F��@Y�-]+��Y�룢�'�ͩp@RO	���>���0ݾɩ���b}BI��.|��M��7T�7k=���=�G!f{x�����¨�e"�_�~D^���&�yiD��=2��cfJ<)<f�I$§?�I�F$%�mr��=��1����xc����!���)����07!ƿ�M��j�a*<e���i.��7��h<"3I2��Udn^Z!H���A�L�0WI=��O���'1�_�Ex{.�-������9_�����t<HHg�Z�Zb(erZ�~>��ei���.c��]����	D��{��<�s���� zF��h�ǯ�损��]ɱ
�y-"��=,�a{?���F���J��0_��ufۄ����������ًLhH�at4!_�,�k�Q9�������
��x���^�������g����Ǿ�����~)���΁�O�B4=>^R�{zG:
��7;I����*Ʉ��?��+�1e��	N����]i�[�i�mEf����-���n�%���)?3�42�*eQ;S�%���H�J�`�c�(��������1^�^�bl&�[`�a-�'���h���kTX�f�~~��*	̼(RK�?�@FLu;7���u�9�͊%�-S�T]����*%)��-[kG��I��!��[�c��4u��\�E�N}]�T	z���9S4��B��:��c�����ɒ��U�/�YFg�:��:�yAz��@#i�we鏟�+��T�T{dzf҉��k�8�f�kL��m�%{E��ʷ�8��w����ц:���}K���7��wF�(��ǺGJ��?��l2����g��|Q�����`�B���Ky,e���x��lb�adL$T�GČ�t���i��m2�HlF$Ď�Yl4l#�c�f�>�3�-����;�w�&�uO��{PĴ��j�VkU}�U��s�����ֺ�ړj�����Ñ�������΍�='%�͙��N�&}��A��T�J���Mݿ>�)�~���9���}��b�����j�*��ԽT-�Qו'�O����̍�<H\F���u�=�<�P������y�M�cf�����ޕ�t�h��8P?B=d>�Y(Z$��_Z�ڬi/![��ljL(��R�0n!~"�X~�&@:�; ���٫k�+�`�[㛄�\���� ��c�����������a�>���A�	/E/�<�٠l;2K�H�/�0���Q9�Ab�}bN��4�3C�^#�p�����(qmߊ�����ĩ���.�wB}��
-�wMW�_��k���q�k�M� �W��a�
�z��9��龸�w�y��jյ���+�~�~�<���	ZZϷ��6�W����I�7to�4�X�Yl"����)Z=å�N�E��|�W�j�![l�o��+�{?�~�(hS8ȴ1T�.n�TT��gN0NVf���\U?l�l�q�x[��6h����o�t��[����]��G�j1�nz�~}8�=>��"��&xM�bw��90#S�����e9Ǩ���O�&K-�#+6��8*�`�k3{����m�)읯;8;k3�Uz9O
|lSo��g�g"�v�kV�^�t�4�5�i~���syt�=~�ϞSZ0��d�zq�qɄ��5-�����u{N�tv0�ո��������c�'�{U�{���k#�"�K����7��O��k6j�6+ά}^�p���p.,��UwbFPUPm:ZY�Mja�RP��h�}�1�N�y2����O>28���0����W����ѹo��גiZC��k���ņ�U~N��#6��I�7Ú�n��eMI�.�7X��Ľ�k�a�JpM0�ir��V���a�v�M�V��Ĝ}˶Kc���i�H�7��L�_B�u�`���ٛ����M7����s�?��.��~��;��
%��z��"C_�~�-�Q��r}ir�us�:e�d��W�5���옼��|"f>575��F����!o����ʝ���Y�Y��Tٮ�E��a����U��d�$�*m	�����3�����z�|Ӹ�ڀ��[V+{�6\wk9�\#r�s�d<b�h�r❟܇�[^����^s���: �г��Jq��5���J�9:@.}־��A�ƍW�֫g���}���[�[dur�I
�-��F[�)Z���X�kT)�B q����A�\#�@/�@H�W���������� Wx����?�a�����S���"p�Z�YY9��:{�tw� 7�\��A "��AQ�~�2j��硧�pv�4�t6���qt�3���0p�h�aF�����]�G��Oa���6-��&b�z*����nV��`N0�8:55����������݁ob��.�\\��ޜ޼��n6\�BBB\`.���������;�_��g+w7;;g'��f�Ξb�����﯉�|������o� ��pqs����n�����v>V��e��s��
>��_���=��}.��=���{j�[�I;;�=��5�ߝ�?��"��/M��f���,�.�����ѯLg� 3��ɨigĿݪ8��>��(�op�U�y�僰���;r���~�[���E͹�[MZ���-�Zv�kvGfeY�d\ݷ���W
�x�%��P%ٷ����_�[ӗ߯
���^}w�~l��:�0��D�o���~K��("M�ߏ$.��d�+��?lT�(*5��[j���+'II�?��4J���n��v�7�G=�s��W�/�(r���Ɵ�� ��>��RW��3���gڐ�'�XJ��9�B/{EvE~�aB��h�	�}�5�]N�*�d(6�aMa��I(�%�Q_q;NTF�:ϩ6zmDDEQs�+�x�Wm]cY~�я�5C�u3r��ß{~�Tg��q���2Fˍ�7�*Ncã3"��\���4���i:-]�Y�{.P���dZ��B�e���X�4D��z��>0��	p�T�<�.2n��Ոx�]]^�̭�����z9]�pO�6�{
�uN3�6}Y=�czD1�e�v]�,�II�.��(��Ct�=��1\d�e�P)���BЉ���ˠ�u��bB�0��H#����@*mg�.A.�R��=��F��_�}=@�ށ f�k#N�*�J��#�:W�F�W<�,�O�d��2����4��ȯ�Ipi������ߏB�G�0��$U28��ei!(��2�L��/�SXe�L�Ŵ�4#�[.��*�E�9�'ݥ�_V�����ڜp�-P	��R�`H1���8�kX<�ЂЏ������L� C=�?�ʙ���.0��.su?���լ7�
V��#�l�߽{�x�1�g��<B'�����4�H�e+/��v�O)�/w�,�{J��jl�cI���<y�Fzج�'[�%�\3]�nI��v�c�8��݋'IZ��/�Lez���f��U�~��ނ��'Pl�!�,V���H�jt�O�z~b��aw�ɗ�'C0a��;�)�n�۫C�R~��p��kܰ�x��XE�	�_�^��]�����V�*�}��V�&����ɨ���4�H���S�n����玵Dy���:�"t�H�����:;{w��ז����8=���5}V�J��O��ʏ	����i��|�����/>W���N��P���6�A�\��|�:,C�A��-���á��A�ݦ$�룡O�ݍ��$/0U��i�K�7 O5��&��LЉO�Ho�g1�ں����}:+D?B�n�~+qp�c����=��@-dI���������L�'��)��;�􉃒�h��L�;��^2^迪?C�9J���;�,����Ĥ)Hb ��E6^f�H|N�"����\��*�[�짚�;���i���co�o�e�0ދ��	_����_b�@�<�RjZ����<�) "!�J�,��>ޮউxsz�Ί-=�Ǘ�Ғ�'�<�p'_;X���(�čw�e2A5:eZXT�]����7h����*�1GtY�lGK�9S�Q�_�9�N�������B�B慈�*K\��8<���ˍ��t�-k��z��P�O��F�3BPK��� 7�<\�f�qP��#[���OH�.��+u�OV��<�VN3�I��(1z�5ǖF�����%�K�K䀈F�BA���\%��w� �!����(\���	0�Y��x�їJ7��ܡ�L��m3��I�Lq+<�Ƙ�If{�5���F�CD �Q���,� �jn���3�[���7x����L�a��i.��D�(&���e�}Í2����,@%�8���`~tz�a8ؕ�����GL2�	8���L��6��5�O�ݱ��G�j��|���y��/q���B�Eqx������UvAK��8��7��>@��������m W6�6Η�yƠ���n�e��}i���ȁL��z���GM:m�52t��tW��6"�z�z濣������J��[܁�L$��UW"���|F�r*,;��&��h�o�`D___�� _a��B3Ζ3��TS�m����1E@�4��8ة���d�~Q#�ƒi�� "�O�:�kyD�e8�NTZ��bQ�o���}���g�{���@�����E�
�EЂ��þ��Ø݉*��t�n.,��f|����|6���ۅɱ���K��sʴ������`z&�r��	�G�"�"���~.�� �숧���4뺛W��dҁEPp���,@��$SX�m܉���� �_͖�Vܸ���9@�>�+!��g�8�2����q )��[|��SJ{����*��J7g�&�~8�9�����4�<�	���Ab�P����J��(Em�;��� �{�O�����D�����t%I[��_��1|h���g,�JM �5�e�ܮ�}:6111����8EO��}U�tg�,hD[w@�4�В��@!"Gl��:�9�w)�>є|��2�t$P�aP��x�6p�f��Xb��ŷ���4�	I	 ��M�L¥�1��HE��
������z0�L�垧����G�4]?�鸢�Ġ�:�58���Ww��ͱ�ui���%VhK���p�L�cM�o���VXx��+�JǛ�/������Z�@A�	"���	<W <������@nDţ����
�~�v�N$&&l�؛bye��:?���m�C6�����?9�GÃ-w� �uN��I��h��rG�a!��)up��)XS��m �_�|��q �S��Д�|�A��M|rh�FK��_�UTT���M��/����gL�=����y���v��98��G�Р/����^�n{)��?�_���1��\Z�������ؽ|Pu�c�����gY�=�k�$�|8�~����(���(<�CD@yS�@Ku'�P%��±_��_�@�C����^g\ԡ�=�{5GH�>5���U����Iq���S 8^�O��}_L�3�e�}��������D���d�^?�/5;"�:QF�~g\�s*�}=�ɂ���o~���@Z�3�}#UzH��;����}�Sc�2#�z�o33�(<��^N{,��xO���,YQ���Q>D�U"o�u�ɹX��OS��?/��N��D��@��� �e�P�d�8u]W�n�j��jJ{'#57��`�z�3$w��6�?����U'B�C6<�fW⢜f�rw	5wn�ƶ�E#�IA�餐k����yљ����{7���臅�O~�����c����M{b�.�
���w@C*��{X���Ock?1w�ۨ��K�Ip(� s�����v�1huoeY*)�2(["�Gt��,�<������B���Cc�ߕ�s�vݖ��˱z��:��Ͳ����\m�u�S�!��S;U�A�դ�"�u'7v�R��i�W�A�!�i�����[V�ĺ�\���J��[ȶpA[�sT�W
�c��d�*!4��#�Oj"����_�Y��G4�D>�K��e+� m?Κi�)>I��I��AmE�R^Y +e���s�Z��MN����YVh�����Î9���Dq �|",��&��㓊W���K/j��ڕ�F��4]X��@�!5��(y�!n�$�м�<du��A�Nسʂ����~fA�T y*���4��1(�秚(���Ŭ(p>HS�-c��{� ��K/-�X�qk��w�֓�:w��;@>���=�A�5&���B]�rWJ�JO�%E�F�\C�N���.{��]^~/JG�W͠};`��n�&��VZu�N׻V^�|*�m�r$�D�q�.=�}�
�{t0{=>�z���%�7ŀ �/�i�W���B�Yvss��>��"��˸�O�P�Wy!g�͹)��C��-���y.�Q-b�����U�ь���t���=b��9��[ة]0�	�z��d�����X���bآ1�jwG�2�=�L[D�ll���օ�1m�p>����mXb��6�K%4j������>`��37"�Sq���e؞�ꨨ���?����%VN�̯u�� �x�V 9 �O8p{ⶄ�=ӘZpՂ�)��X�KXC�ӽ�*������/���f���;��k�w5������H�l%��Oaw�@������@ݠX�rQ��ƕju�E�����^$��M0��2���yREq��rsh|^x5��X3nO��+�V~�׸�I���ק13���
�4�f�g�����zX��U���:R�}�E����U��;�I>��3��9C����9&J�L�`��O0�>��.�w�mbJ��,,%��H��cYD�]G�,�y�C�p�&=Us^R~�h�R�kՖ'ˮ_o�00T��*8�ೣ%(�1qF7+>cq��V[����&~{�DJ.+�>5�W��cּ[����t'�G�{��q��w;L^(�I�ʂ�9��s!�p�b��c��(ܮ�����aC8X����Q��to������S��e������Y��*:3��f���Q��_l�u-$G�Ec�� ����Ji!���U6}'~@����bx7�����n�O�~���a�WPC5z��$�&�L��0��h��rG9�2���3���e��.q�� >9�f�<X��mU�Q��
!\�3[$���
��C�_e=i�)��� F���)d�.������Q����ٸ�>�ëa�R�l:�?�n�YKw(���~Q���{V0��]����ɇ��C�6�>��	��V�Z�e�λ�r�������ix;}i����"Z�?����V��`��4��\h���~�
��k ��۪�*P;��m���$[�f+���f���a�?�ߝ�������^�e��Y�?j}�@����i�*4�����|J?�*�?��d��,��A~�䷞�������]�3�'OF��.O�H'��x8U���u!	���'��M��^0����nD���?#�+L�b��W�K0fsxQx���p)��˧�{�Co�hH��Q���gh�v�Yȍ��-q�* �8���)\�0�X^���H�|�x:��f~�t�V(����[;	���� y�s ������9�lo�sx�5���Q�ar3zAA-�ZOC[%��c�	�`�$R9�D��AV_&�E}y~*�(�[��Ņ�甆�Ka�}8�!���(�7߭�.�7;������o\j)�Z�i!>�{�M2-K�lBPgϢ�Ņ��
7�R%�?bGo��q�RdJ�g�j��u�:*t]ljI�i�@!��(:�>�p�u"���~��p��^!���&"@��Q��Gʍ3����Q��(s� ����m�j�{��zAv�uO�Q7W뙕��Q�P�`V܏�C���y�;$%���[)Oz�̐x_�yvϣ�»Ȍ/�ۣ�����6r�~�R��EfXvK����Sv�=5�a_G*L����pN~�$${�L�3+�x�I:7�˩��yu'����~��|�A��y#Z&a=�� }���9��-̐T�d÷\$ P4 õ� ��7@�����V�q�&�~�����S�e~�۾v_����8�T�0�i(>Χ�����B� Y�r?m���C#8�OU��u�e�A_kI<�`�R�-|���*@R� *؜2�r�CTF�Kb�EH�r�b� C��W:��BH'X{m�r������zS�#��L����a��VU� �gF��UW�����YB52��I����$����&����z�黀^�CZx󕁐ܣøSkG%�u��[�9C������8S���+�V
ס�Kt�m7��k]��5��i��e�w�B�g!.�ZO<|�G�:�8�a|��q`�2Hc��!�2�P�S���diIY��3�2��܈*c���'��?����P*��z.u�4j:|w����\|��u�Ζu�]�>&�����V���Q����������	�M�7��)�� ���� ��lfx�jl�a��o,��G.�����e�a����=��y��o+RYPI� ��6b��
>'?R�칯�}!���Ġ�]�L�vc�%+Xm�3G�Q�~^:�� �ŀJ�(��Q���۔H�0�B��q��C���;���������#化�L�Eo����-<9�-�R���%��ȱ�`���$EI���bH/o�i(�Ǝ�Qj����У�L�M#���cqx������3�υR%}=����xYT�\���o�O֜��r�?��$�½��5q�(�j����cf@j���/��$ӵ��/��0��d���H;d��XĮћ#���"�
�#qg�v�
�7��.��#�3/��˳^S�Y�i-,;M��5�)��V��GA��Xe�U�.�ٙ�γ�+++��:r!b�����2��dɘIx��G��D���R�/�?C��i�̊#�{�ɆO�uz�r�҇���o��ό1�>!%Q����
��1���'aڏ�x�m><����e����;�d/J�٨t�������=��z�c���ڠ2W~�v�&���ef�P��;U��C��"xQ�Z UVPp�6�*L]�򆽃W�(����u98(X���x�
�����<lD�:7֗���S��ŀ����	,CVq�? �;�Hf�O3nJ�U�����j�Q� ko�6b@��uM�4w�����{��1@|��������c7��L~�x��L`�n�ϣ�RL��_a�1 b�GFMC֧�Cyt�'��Gs2s����Gۺ�Q�^$�C5o�M��&0��'��4څ�I���l
�l��5B���+A��P�N^�'�359�8�<�i����u�}S�ܣS|��9M��XY���<K��Z����8��fTKh'^���s�Ok4n�B�p�9l��V�d>/�����C�SLV��Y�iKI�e��m��ա=Vk)��]��;ۉ�u���3���\<f]�pS����u&˟a#��7�4����[��A�M�OM"V�Lk���.�$��ZD?��;��n�^������;�&���+N�h�Q,_x�3�=��T�ە�l�>�P�=�67s������hŶ,�b�+�/ױ_�����@�����]�Rq`��Z�p 
3eE�M�Nb]�,h�8���N�0?;�������2����l��L�kzW��Qå�|E�l�i��d,��X̑���O>��x�(M{9�[ޞf��;��h+������$�N��X	���-��(���9w#̆
�0<{��o3��C���}�q�>vRS�mL��c3�(ԇ����|��wE����G�O/�9��JJ��#��Rw߽��)��;;�F�)R����Oߔ�i�����k��)�4�����'��Y��Q�AN�M�O����W�,��y�[Uo�n�?>�
�����C�/+�����T�:C�6_�&]ӑ�`�
0r�����J-��I�tF��4��~m�&��B{���XD��&R�9��v8��%X�G�?���X�Y�,1��
�s�X,X�Q�!v�����<�#��6���*�yA�яx�������؛�o��<��銊�HU	u(�C<�b���K�ˉ9#TQmj����?�8�#L�'�L�2K���*���6�G0�#��!A�����-�uh��c]����k�W�A�m��$�9%��Wt�|ֿ|���|k\����"���jQ8تa���"ng�Gt�Ϫ�V2�=��+���b��t�������OuWi��IV���N���U&����ߍk�Uf��^ֿ&�c���͹��oKQ�^�:ir%�r�1,�� [O�+tuǋ���]:����]�ܨh��/�<"OW
�zϼw;-��k���F����8B�d��;w�4����eI���i߮����1�u�rX�����7ۂ
sa����u��a���
L��6^7�9;[���(�U���S�Hx�趩I�-��v����@���46�67�"��5���j��~�³.	�2���`�#]e��3*�˴Y��F��v�p�\����+��׬_�r�������0�!��k�v\n��=M��cz�[N�H_��nP̚Y�V&��]�ȷ �������Q�OG�.�Y��O���ਝt���o�����SU,�T/���a����0:;��@�s�u���ϻ�
9ڿh���%B��PՏ׊b`����:TT�g�y�_�����H��疩��U�������5
�����p&z2�%�a�O�U�Lr)D?����pq-�jI��2/RCbވw��Q	��N|���	��d��p���R��-�.o�������/PF�@g|��J��t�!�[=|dʉ��#��9r�wv��"��ҧ_�w!W΄�Թ�Gz4|JN��;�=ھY+]'܏�Â�i�)`#n��9�`k���R�K�\��,T�r�v�dRSn��1���X(����Qܳi�|��tX �g׊*TL�Px�mu��&!&�%�������e�M�y�~��<�&��z�3�w�+��!��a�=�3zW�>���9%.��TLw����B�׀��Ə�*��D��q$�1D{�.*�?�e�9�p����U)�yp��	֦#��I��۫�~s�:t�9�C��.��V,�s��>	������ZѾf(gɞ��o_H�{���Pe���Ȅ�D|���ÁͿ��9{	
_�`����ۖLvH�J�dUy��Y6���P�Q������k4(g�
��A����S�VKY[vB�t�hp1����2��A�O��!h���Ϸ�&a����Z���yU쥘�Y����8܄�Jo�M�n�K�5We�J�mKS��+�#�рH��z@O�Ep^��]-ڱ���4Gen�v`�an�K=�h,[����?��i�ju��`�s+�������i�ئC�Au��8��)`9�,B�h���z�&;��ELnG��(y�c�Bxu�����Jq>g:� 0�ĤYk��0K5Մ��|�Ӆ�z���F�f������V������hg���J�m"k���!�ņ�md�4�p��^A�
��R��m/���mSC�_+qYB��g�"���Si��F�D֬��l�����dy[ߏo�&7���}f�TҺ�(>�*������6.;�[L0�Z��iE�=���2�8Uߌl���׻oZ4ʱ�%��������Dԇ��A	׊ޕkB*�U�e9lj�ޛph��x�����G�Y4!��f����9�8�|�d�e��S�C�x��F��E������=�zv�Ո�
m<"ذ��C��$f�pL�	��F��'�ЗM�W��
����
I��z_濕�� �^����9|mߞ���gR�2�B�v�%�m��g��@:U��b"캧זv� V�z!U8u� �)��d�0�a��+FH`�ApI)�Bb�!9\��?唝1��Tba�>�,u�?+�RS4��u�,�Sn������AB��"2p���cZ��̗�~T#8$�� �\�[a,����~އ��c��R�$%UAp�ޕ�L"���.���Q��%��T�,z�Ua��o~��Be�}�5������}s������>G=�^哈��91���ZiF��!*F�-��q����l�\��
�\�@=ݻ����Q�Ħ�q��0�����>6���2���\%m����^a�{s.o�=W$�b�(�n}���V��W�m�q�_,&�6+VB���f��ڸ�`���<uV2����'=X�X����~��ᖒ��7�O7��V�J0���>�1���]O����e�6:�<�K2Gh��^T���5���d�c�Uu|ᗔ���La��ȱ��R��tc��,�_+�.�?a�ϖ�wA]��o�55�k���B�=��b�P�%�Qv��Cx�G�_D�t���&n���_Г�i�Ǜ�e|��2���,�/15�fw)����R�k%���d��:0�	�`�z�]�3���h���ߵL_�6f�}ں��6�nI� |�-?��ļ���q���Y��`���E���E��?�3.�ܯ;c�;,��v�Cw���q&��+l4��ws?��j'���2�nn�y� ���l��yk�Zm�@�=�]4Nss'.We'Q"8�X~3s��<�{�iL�L��r+0����H�jȝ������G��x��P�n�rp�@�1��u�3F�5%|x����ċ;�)�#����Q�}v��O��{Ö����B���"�k��a��� �Þ��=M;@�r�>���_�Q.�ă����{��Le�;�R���,[������1��ү��r�c��hx���'�?��ʛ�_�k_�Tǃȹ9S��ٽ:פϫ�3|�b��a`+�/����ӝ��nI��)bF;�vg�k�:Ѧ�py2�>q/��T����S�ͺnވ<�:8���n�~SE��6G4�ܩ��-��Dj�-�����C�^��(�0��r,�gi��xp����M؊�9(���6>��2E�A���d���C�'�70o���r#�7�2[�A�ٝ����K��/ٓ����5�7�c��ǫ���?oI�n��qh�c�jS�u�QK W����嗀8X���3O׽:�.l�\GL������j6�f��QD���2��W����?�݇,x���������	��uC�*6�7'�T'���z�x�x�A���%���>��i_�}c�ޮFE�"r�(:���9
��� �-lO1�m��2I���|��y�6@�^R*�xe������o9��(�xUș��1 �v��5���-d▛��5�W�o��N_���!ۣ����Dѡ'������ǝ��~N�{wr�	���Zt��۰�W�3���"���%EY�~����}�>��_�4t�zbo��	_�A5~�x=������������~˿ft�韻N��D���p�ӟ��2�E�����s�K
9 �HC�PT����fx�|��Ւr�]�e��ù'y�r���x��@�����rѮ���K��#��]�|��w�u�t�a[�N7Snu��r���*- �����ա�s	:��g���91ea-��(p��خ��{�H��� �N�R!R�	Fk������X��8U�ЄlN�Ьk�[�4�5�Y��T��F�#@�U��G(�����OWݴ�!���r��s%xy���WX[X�+\;���4ҳ�R6D\�*��)��С&�?��*}�o4ߋ��ͮ�N�a�_������|�=?�?��ǁ�f�r��oY�	}>-DH%�B1+q��Q��չ��qY���ɔ8���-z��~A~��E��{�}i	�Ve�#�,�M����������ۙ)�P��Y�p���N�?����˺��D��O�z	a㭧�X���yʌ�؞Kt?EJ�Ȉ��ş�ܳ�7p��=�н*�s�~}�ٱo&y�,�ȣ�qE� "�%+xr�i��̕R��-qO6�]���GiG�fv�:Z1<�p��	:˼䐀BEذ�H�h��&�m��eC�4�vq�%3��YWA���q4<�Av5�<J�x���v��{�������9�z(j�ݜ�wY�8χrS��a���.��;��h�/'K_��!��f��`�^,w�����+ǫr��zs��U���2i�`��hB�U1W�Q�ݳ���Q�$:|�@q���
H�\	e����xl-x�am���́���D9~{��3��е�]�m�+A�LCHcޏL�_O�'��$�$��aG2*}� ��
�-���}akD@�z���� i4��4�I��
�}A!5퐜�W��Kx��**4�r����i�-f���!�Dv[�րE��]���	��ȃVj�+:8���*ॢh���l}1�ޅ���I���~���۷p����cyL�����6Т��Dr�.+Q08B�6(X�G�m/}$�v�lOk�r�U0� �MJ�1ܮ�~R#�֘����k�z�5]J�g�+6��*��:Q�Ë�lz���.�����~�9�O�D�,/s��e�כ�r�Ɯ��J�>�?Ƃ�4Gd�o���H�>>2_*��S�;�m���%RX�U~�㙔<�A#z֜�� �6V1H��{a��k8W"�N$Wۥ{!>� b�Q�R��Bs�䖹N��{�d{�@B�`�O9��I͖���͵556^��,�:���X|���6���am��<T�S?���i��N�r�Wc��X8Q�X�(H��z���M�v%`�g���F����C�������ѽ'�80��϶:�;,�-�Ǆ�?>~-Tۥ���6M�sP�п)J�l/����Vp���6ɃB}�_����(��'��ө!c�\~R)��C���F*3�YY�����AY��(������p>���/���ݱ�.�5ެ�q���#�Rs1�"���e�t�n|xC,,��MI"~�g�9b@�S  ��u�吕(@\�����%`�*{(�� ����a�olP���4r�����F�#���c!�7�?��x
�� ٶ���X*�U2��o� �!���w��쎩�{Ìv�p�+K�������2�70���
��!���B���A�J� ��*�$=�����BF��w���=�Ѥmqӱ?'T��.��]�`	��L��e�dN��Q|c�ͨ�O~/����JK�����E�-��c������Q�m���^�˭c_�
��擪�����$�M}1���[����}~66eVVV�V���T�V^
�@)�~h�������Od��*�Z�Dߪ�(=NH��_�naՏE�����"d<mIPh��̓�-�8��h0"�������`�3쐝KZIp�3�4jd`$�z�7�����з��g��2��Կ��BnAk-\�HP�����h�묻��}��rݝ51�	nh>ˤ¸uq/��>�Kꊝ� ��5ȶt��tLq�&dP-a��j����r�w�������L0��
[G����~�m�O�0�'q�6�T��_�IߛN�%���p�/����Z���/L�n�d�J���Ĵ9ė���b�R%���(FX���S���B8^V+ݖlv��H�4)�t(w��ч�8�ї;VM���ea�𝪰L��o�*��a���ʒ]m�*�#{,Xk��%�̬u�]����pJH�}��I�ueQ=��)}��X��.Hn���]t�?���I;U^~��dL#�7Q�1�xۏ�:͏�i	�J���
�g����l��Tz0p�,�k�B)P�x��$��r���|�kE`#a���V�I��ù��,�g3��_X<"*4��<~�ٍ}#?i����[��W�0���7=�^l�
�Mk7ă����Qa$~��u��憎�;��opQ��"_� ��GO�C>NfJ�u&udԝ�؎7�8�m&l*'��E��T�����p�n��Oy��'a񍁊���[�K��q�6�K��7���uB���v�W��HC�2��h8�E���\�$߆Y�J<6��	�	f;�La�]Q����ަ�t/��oW�;��{ci$���rq�`k%z>���\�WW�l��	�l��YO�-�V��x	����(#~9�<K��H�i�����vm<d��H�
���z��M���P�����s��yn�[�+9;�:��R�[�}$���^�\U��	��7��p^�~�^��eSgv�_�e���Ø֮t ���?қ;���M]3��;Wr�O#�F-f�$ӑ�~���~sX��7�y��l��M.��|.>o3�3���t��oM.]԰"("�#��4E�MzE@z�]JUJ�#H�ދ�P�wQ:D:�I ����{�s�<����/p]d�={���ړd�������H�5YP��g>��y~�4r��N�n}fhq�H��L{�19�&Q�G��`� ��+���J��p3s����8�p�ɾ�(H�tϱIJm�J�#��Dz�4�:��dd��S�V���/1>c�:�j�����&�6g݁n��Ƿjv'��y�4��:�ƨ�d�~ ��.W�ցm1�I�ዶi����1y���o4�Vz���G*|8�C՜򹡾t��5fo9d���/�cǮ-���wo�<|���y�-5=���
�r��>ދ�� ���Jf�ٌp!��ª*������V��}P����#+y�<��5]]c>����ɢIW$o����"�k�5�%S��F�[;�_w~^*�sGۭ���̻B�.v���lL��'��$u�����Xm���G�V��p����znX����H-��p�nP�ca��%�4��Q%e�g�,�����7����&s�Zs�d�V/���g𬭬=�Y��	�(�bR�U����]�X�T���F�xt���\b��N@�Ն �ݗ;F�$!�����]:nç66y<�������4����X�V���!��:W�`�BqI��$us,�^��S���������?�|G5�~-��a�F�y�E�߮Tþ?%�V�LvF�Vs��ߠ.�HQ�C�+�SH�6��,�1%0H�+�ul�U����}�ͭ˰ٓ����|EA��'&-�.���`�R83������k�<-�:�V��׫��q<���e�i ���Ո+O�`=[<�N8�u��=_z�o��=���H��ޯ�K�⪗�A��8)z�7�L��N��b���@�(������|���l|��IBJ�]g&R���
-~-pTq��{F�~l�Pl9���+/婢�M�uQUӞ�L�{�¢.�&�(<"ԥp-';a+�ѳS��
z��?�%++���?�n&L�s۽8�bH�|�3���ME�,a+�EϜZ�i�J���6v�a�ٱl@���h'�Ů��+gT����@�\n���sBAn���o5jP��,�N�q�em�G-��9$q��eև���y݃)�=U�4��v�j8�{bi��K��C�Co��KkG]���O�Z�w[��e�))�.��I�ceMo�8�@��]�ݗ�Lj�1�摮��(�����~q����	YJe'��ͻf��3/��x����֮N�8�9J�4��$��Ȧpg'j�1d�oE-�sb�oa��Øt٩����5p�V�=m���7	D�������I�w�����ԋ��O��<�K�lC�K�M;}܅ D������n�`s���G&u�I�f�e^r�����G�_��Ρ�S*������م<�!���b2�8ۣ����'�$��;��w�br���-��Ջ�K�X�����YYq�<�EP~)r�P&��'����c�_ߤ�f�.m��Mv�l���Q�㊡��]��J�|Ti��q���@S+��h�p��UF+/T�����_��Y?/�a��֦X3K�� UG�k��d!O����`��O5�k.f��Q��mR�S�+n��J�����8e��5�����a�Kn��>�����A��J߻���yۇ���3�V?��Y#�Ԡ����w�DV���(OG��N��'�MҬ�P-i5��gwqȴ�49��M3�pEe���MX�^%:�  u9� ����dv�yn��On��B�8��X�L�X�٪�\�˞��ђ��q�K��	@��b��7�ʹǴ�vj2Y����;	�R���H���DkG�oDQ��C�R��L�8� ��.-���s��$�Y}��C���(zw4N�J>��{ݨ� �]'��ix����U��m4��>\lz�J�>{ȧ���o�Kp��#n[4�Z����G��|X�B�:ѯe�Ӑ�e�_�6r�FTv0�]�ZQ@\�:��f ��J2A���m~	�
�0ވ�����|1�Ɉ��e�~���z�M8���y�������(�ڬ�Ӽ��שD� u�~3*<h��@]� A�X�֠��7K���KQ~�0���	�Ԫ�M��-�#x%�P�L^���@�X� ]N�k_�������:^�z;�;�9-�>_br���#��C
G���:�3�xBw�C�{�i�lE����Uu������w6�>}
�`��9�!^�K��?:�u�t��Jg�3�&t<��hR��������\�B���p��y�����I��@a���@>���x=��M����܏_��j3J��ȻD�b����7fOt���v���L0>�&yN�W��^�F���\�C�\��$(�ui� 7 ���Y�y�Zy{�i�ɮ�~R�̥L�(�~���'%��w�{N~��v��;E_����`׽�#�9�y^�t�(�V����*��0���Z���jTs�`݇�G��e%4�SD�I���N�R��;y@�kh��v��U�����^w������"�Tr܊�f3��2n��^0������T��CLsC9L	Kf�֬���5�@(�z1�j���ON��%, p���>�鞫�ʙ���K�m�T�ˆ��������A�w�%#~v�R���>�;=z�T�� Ք�"�=d,_�+*���Nނ�^�!'{�u8,2/��X���+�r,n^�UoA�n3ܤ(�B�D�W�%�� �^Ķ\)aML9��g:
H�_�0����1����#64[MkL��^�G��=E<�Z��xw	���O[��ޘ�blJ��K���|�4���bm��	��I�)���&�~���/H��|�����<H��w��;�׳������*�,?��ci�y+����1@}H�:���y,=�=��E�B��T�v��>��o�d����9��R��˳�FwA��"��� �����1RֱWX�)$����E�*���?(zI�׶KѴzm��k[�'�*)�����|&���C0��&��?���d���:��37��t5����=}��n(��r�ۃ�!���"窓�ջ�T�Zp���_B���wT(E�6Ȼ��%-R�5�y�q\K��wB)q$�ݢ���j���Zy�[�âa�TO���5�r�w���{MmWR���N���rxaƻ�u��2z�rohQ�����V��&�͔d���w�8���T�� �⏍�E��H5r�nh:Ͼg��P�åZ��9�Lk<%,�6�a��)pҮ�@����s����}�-@�g���Un1"U ���Mh������e����s�ں9x ̲z�V+���O$*e|a�U���/((��?��Ժ���۫��<5戓�J��{#\��ak�.�}д���g�|�Ua�^=��&��F���)c���I�3�������ӓ%w��,C����gǘk�6�噳�{���6G(˒8��h&]�iT=ԏ�OE�`�T���T�r�H��	3ػ�)�M�D�C����R�����N�)[0 �M��%�e�.��F���RN>�<�Lu�Ya���X������o���d@�ւ�Us/��R� ����l߭i�Ն�S~�c\W�~$2���󟎌�7B�P��g^���߲���P��$E���-B��K^40u̑��T�飭;��S��h����ʀ��mz;�+���$���wS��
Ϳ=�;Wx	S[�a�y��tް�����V<�+I��d�<hU5��9���&��]�V������?mZ�1
X���C5��G2���G�Z9�+�<�D������<������&��1��
%8Fc������Nƙ����!�a�.�x~��^�}��[�9x�5z�ǗL#*����h��E��9��KI#﵎Vn�j>*���>տ
�qk7]�iyTOK���| t��VYw�ϤX#C��u��ȀZ��9���V��!:�	��k9j��e����o4�Y�8�4� �{�H����Bi�prU��:�fg^D
��(�f�ky5|c�S��Df!��G��}���9	u�� #Ĩ|�]�b�.~ /K�b��*����N/�v���\ڀn�C�6D�0߈W�&�m���ֈ��%��������-/������z�	y����w�`�͛��^��Ԉ��>d��-�b�Wb�W��Lj˼�`�h�	i�^�Tyw��Qβ$9�M�q�NnЪ~*o;5��6���g�2���Bp?X��|[�6�:��U݋�i|W �U%��<2����O��V
C<WG�亃����<�~	M�-�,��-��D��hgJ��� T�5��>���T��LG4�%��_ξ%��K�1*d�kȒz�02	�*߱Hf�:��<h�̓t�V����;��`���{>�X���4qb�MY����`g)'�
�G�N%�;) ��,���${�ˠ���]�'�?O��c]׷��}���v��Y�h��0_6�X�X/qUJ]�v�ɿ')<_ơ���ꐬ'��N���o=��П۶5.�~ĳ�@JsVM�ǯ��6�IF���Əae��*l�:��US�P?��o���;�u;d:Fϳ���JMfw��h�q�O�DI�Ƽ�p��������[f9��P�@����,�Uֵ݁���P�3!(0[�^?Y���zH�Rݧ*���j��$�z�5F� ��)
v�Wdt#!�s�=Q��8؜�Y�B��[ {S@G��~���i>�f�J������`;�e��޺�����~��T@�k�wQ�'��O��t�hS�Y^���<o����Η�硑I�E,T��'�-�.�:��q�z�s�e�页Fzq]��z�Y h ݰ}K2�������ǭ���C� +m�����Y�cu��/<��]/I�����Rf�_P��$�f�{O,O@����kj$3�Z+R�{p���������44p�
h�9��`ӳ1'v�+a	�U�N���� �9`,��Ee�p꺓�l�V�.	q4�һ=��߿�:F_^{�ة��'!3(�	޷2��{��9��y��c�?��w�/# q��X�,��ux>�4*�r2@��!�W2�^��;m�՜�<=�[mT�ʞ
[MA;YzL�2?��\���;U Z�x�(Ј[f-�;y>-~-K����Sr��7�b$<�9Q"���{��0��I�;@n�3ʽ2���JV�;�Od[�,���-�d�O�'��z�s���΍�{ؖ�{�^f�2an[ۺ�|���r(Xd�b-�q���'�x	�"*b��2�����lEW^S��z��+�%9�_����{Vϳ�c��i����7�w��j#����S��{t���`�X
L#㰱n�)��цxn�OAB�r��k|
>�5�x��
��9�K�O@1>z�[�Q�(�~	��s$�o4rtI~?�/���=HQ�9rRs��m3���W$]���k0���˹U����K��f�<K	)R��[��)��Zό,ݏ�j���Dg��ǥ�W�/�l�1*}��,t���3���\W~�h�p����w9�zY��P�ab���c��뤿g�$Q�ON�U�kp������s���=P��[οM�I<9��3���?˭��T�T��cR([\0X�	C����@9<)*�j�NzT�w��D,f0�o��Eo�� 
����m�B���v�Z�i���\���ɛ��!NE�V��Ƥ`+�Vuoa�ĪW��`&s�O��{V�%��{��C�6�s^\�O���0�%/����`��-Cߋ�?�n�=�ҔC��OxU�Qc��'�wE;�&�"��j?Uu���
�إX5gxQ���g��&-�묯�C��{�F%��Vb�z���KkL<!���~�`g������!�u���8��^6��s�.|4�]�;@��2�U�S0}� �����>��O�F���<9 z��/��_���m]J֝4�RSٮ"b1�/�Pt٣^�5�-�)�I�;�g�6M�Y�ԵUv��a�^#;y�V�����9
)� ~ t�;/�G��tMN�|��VG����[p���2����4"�XS����jk�~OmK�+ >�';��N8�"(a��[ʙ��D�W�ҩ�+�^�JA�𧽿�>ue�U+�h~�����<��
����1��"�F�W���� W��8܏b��n����P��P���ܛI/���]3������'L��k���*�]��pϺ�N���6�h&�]��lN,�,OX(���)�
��4�Xd޶���c�`V�{�V����Z �w��B���vڠ����_s=v�,T��#�� d�\�1�h.�LRt<�Zg-H��X���-��� �X�Tm���P#�<�
�v�y*�ς���$�D
n��B��H�Y��"Ցc��U�O� �p'=nEȖ%����ۯ#���S����e���V��Z�\�B͈���R���eaǽ�I;��/���w��!�䑟�k��Ȃ��4��iJ�*y������1���KkӰ��g�I���@�#ו�^A���"����E�;����e�+����(�R����s$�@��;��N��t�s/�L�Ahq�D!�V���e\U���t���h$�!$�y��ۛ���+��r�LF���=��n���y$0�νJJ�/NZ�y���
)�W���*?:0��R��E�߸$:�I�e�?>A��9�6������?�-�gж ǈ{.�N�(��$-���?������=�C�g畫�zlV�לO�%R	II�uZ�:$gkƓ��ѽKH�m��%+%e��������l��UZF����N�:�����3ۯ�_�~�Z�E��̌V�;;O6�������{�烙M��L��'��v���3��������Z����bF��MC�	lv�e�[r˴�q
o竮��"K*	s�Q����e���S�z��k�|�L��U���nЋ[���3,3Mk{F��<�e�1D��Zڽ6Ũ�6��E~��!D�A����`�q�ݛL�M�
��?N���5�f?Ы�T�c�R���E]���|wW��JBJ���u�����é�+�S�=�dI��X���$��}~u���pJ�{�'�9VU�g��%	�D�8G�f˭o�t�7��9Y��r�=W�l�f{:�'I�˨�<���Fg�=i��_E�5<��T�2B)�v/�b�Fڟ�<�t>p�x[�A�i�)�e�^,��0_��%<1�8�>!l���̰����O�I�W��:��j�b�p`� ��F�y��_;��̊qAǇ��p|"%i\�ɞ�ͬ�zK}ww���R��uf����=Lj�k����C�b�4�&�n�M��Yce����
ԵZ��F�s9�6E����^#����$�H	�@U����eL�1�����ح��><X����g�3%`r���y]_O��*�$�/u}�[:��%�kV�i)F�ڞ���~
�ш1�a���9����::�U�7����T!פơ��U���떽S1��5]�0c��-ޢ�ag�kC�N�_�,�Dkh��&�_Dn��Z�M�� %����b^���ǚ�y���wm0�[�1��0��-�ߗ�����o�$�K��,��_���+�U����$gJ��M_��Z����;Hг-K}�V�T�~����b��1Im��!�
��z�����-�xg�ZN0_SS���3��U.^&���˿����򳓛�&6��^=S���<d�RC�i|A�߅\���|��0�Wj Rz{�.t��4���hW<p��-��N<2���r'Ƹ��3�5�L7��(���{oN،�mL�2�T�F`���}���NAY��gKK��-Ly���WѺ�b����.�a�i�C�������������t���G�<?2�qKD��eZ��+�1�f���^��źǄ=���H:CH�?j7�
o�Mw�#���}wz��0���*@���;éj�.s���Q�󭜖n1�� �:��$H�nV�h�@���̟��}�^���} �a��K���%�|�$�x�Yn�������8��@��j�tI��Y�=l~���,)���d�Xqę[�I�����[A��.�Wb�TL$����ѽ�~��/l������<���<?�J����cQ��Mr*dH��dT���ˇ�\�C������̮�O�4r<)�i�o&�<AZ�W
B�ˋhFr�#����n��m&�)����"��  ��X���H��~%dc�:��OK����)��C�ޞŠ�`���C٢~�/��4C6��hM$
�K��;�Q���*��*����&K�P����;�*��b`��!�~�� �l�Ce��ܿ�ȝ"{�Ӈ�
��5娪 ��£O%��D}�=��Z��%�9/Q-[���Ͼ�7�Iu2'��b���n�v����'��ʥA0X���%�C兾 �d����b,3}WӪǸRBOS�oȸ��;+�'�ȷԷ��~X�n���g_#����`�ĉa��kӓ��RI`뭴����x�h�󃖝4Z�W�.����)���Tm��7�	`ؕ�Dr�|�tm�~aߍ:x�6�ҝ�~g?h��~�/I�|�3?���L���Tٲ��X;��?Ҭ�
��g�X����C�%/c\c���v��[���z�=h�НU�#�s1���!
�%��u���8��;���<<=�-{N����'g|o�ѬD�m7�ֆ��8�M���G)wc��7v[�4�-����3@U����.�T���hْM�l8ƣ��6o|�[�7JeR1�	�C�`8����!>�;����^�	+5�i�L�;J��U3c��?�Cً\S��&d��+nL)m��>�XQ�d�������|��K�� E� ������Y"N�}B��?ԣ��f��(#��Ҝ�8�Z3Nk��		Z�&1�;O�2��K*�6�SѺ�~T���V:'������W��v+@h��Z\�ǞPm�=�.gߗ��<o�O�?���8����tA�Bk�m�(7�C���)���y�w�b�� �pB��oq�='�s�v�G��DY�XA٨qi5)�����a���\R.��ulF8ӜI^�o��W���
=׆��J�u�Ȑ/PJ�L��O�/�!j����	��B��G�lN@lʝႱ��]$�#|θNK�EY��z����=�S��m�r�%6�L"���Uq�6�Xrk���eͧ�]̨��Qv��7�s1a�W�\��9K��G�̉r>��k)
\�f�^|��e���"�y���~j��.�c�~
���JRNJ�Y���˚�ƕ�XY�䳲��/7���d��g�G��F#��u*�@@����ZF2�@Ʈ�;�
���|�M���慝2 (���p����uV���v �x��O<�,I+�=���
P�o+����f�!Jm�Q��D=���ӓ}HsD6��6�f��C\	��e��3P���9��i�LB�l� �%u��HЭ7'�g�4�to���0Ycj��D�)�6��Q��kj_��R(���C�Y䤀�h�Tz���_n]�=��јs��3�\g2���&�c���WA����������u��PK   ���XB.7# � /   images/1d5cef6f-7e1d-4016-8cd4-58d2b051ad75.png @翉PNG

   IHDR  m   �   ��l   	pHYs  �  ��+  ��IDATx����de�6��P9tW��Ɂ	��8d$(�"(���V����ak ׸`B	$�arΝSu�[������]����ί��+�z����9ω�]x�W��Gw�W���[����"�y�cA�~��gp���b�6����a�3�/E&D\�G�������^G?W/��]�%K������&}��w������_��ۀO�s��Ȩ�L��z���r�غ}�J���>Rqm���:8�D$��B�Z����h4	����,�W�TE�Z��JpxQ~��je�� ��˗`|��U'�F�Z9��^�z���;�?�nށ���,6o��q]���q��ÖMULf�hoI�˟���o�חى�.?.����>y�IxϹ_���9�4}\q�B̙ӄ�4�͹��=/��cĳ/m�ן_��;k���\��RQ��DC\�j��ێ��I}>��D�F"�
��W�ڵ	��l�E�+"�����\�g�G����wT
�YC��|ݷQ!Y�,��q]JY.��p<�0ŷ�rg>����{�VC�\ASSc�YT=�H^)�j���
��s��L,E]&��W�~	D"a�exUsm�be��m����qr���qxu$Q-N�ց�1}��	�2�ۚP����{w`v��(WmMm��
�n>�rB3��HY���~���1�uء0e5�T27d�����S�J=שS�}�C�P��ͦ���#x��T�ٯQ����D\��:�S�$���O�vl���m�Y��ka�v�(�v�φ������y>+�r?s��F&�P�2e��ox��P�{���D��4��8a����a�~�c(,���5~/�d9-���^�s?	׏��&G̚Λk�����4�h���r}�s�F��Yi�
%lX���F��S���/�'i~GB�Ü�x$�j�#�[:�Q�^�|;����/̉���,3�in�J�r�#���9?u�
�?��Jͬ���R��jus��X3�5g�OZ��q����q'v�>9�sX�݃T�Ƭ�6L拊�^]�˜w<;�8�x/RMq45����|D�:�u8��j9��{�����ِ�����	�P?��X4)�;���ⓟ:�73f�|p~��'���͸���c��s�pڻ���MR�]�s����\��O��@�E�3x��>\u�p�~�.��r/>|٩H�èA6U/���裎��[ny�vn��`�t�b?q7�c�8��s�ӑ�ց	.X�H\7�l�Z�N��&0��֫
�ÿy��J	��L�����;�B��5i�[y)h�p��??w��:W���<'���DS�R����!��Z3gS�:����Ps�X�
��������'ቇ�������_��:pV����e�u��~�Ϲ�p�=o�;_;?4������B��G(�E*���e`,�ja�q/Fs���yp�"/���"V+�7)�$oF�s�f��Q�J�T���2��7}1ƍ\w!SW�v�3�\@&����0�G!7	/�N�A��!K N�P�A�\U@�f ��q�
���=C�1-��d�lV'�f#�" M�8�(sS�ON�1�?�k�Q1��O($��D��9G#�D�p[`��שWcw�0?p�Gt��5C�U��a�!A;Xܨ>�N%V��l*���+�|.�M�!�D�	�(�D�5� ����a�,Y:+�a��~Հ��
(��FuQ][琊�"��u�	P��u��s���8�:k��*�?S�7)p{\�J�D(�{�<	̖-D�5
��u	T,��(�0+�]��[���0:����V��y<�KEB)I4��*K�މ� ����3�����G�@��y���n��[�e�6<�����8��}M�s<���麟�(P���\���9��F���T��'l�נ�*�B3I@��5ʑ��Z�Î�º
���S��UU1Z�[�5��NA1�3(Ն(w� �n�D�
'�C�781L�L�հb�a���v�ݰyj�������C����P(P��('MȖ�!���X���k�l�)��a�wc�A�v���'��7o��w=��?��}�Ԝv*�����/?�_'*�����d�!�����n�r�X�m�=�s�9M]@&lڰ7�|'�p>���q��G��g��������	_u�J|�{?������=�0�h$���n�a���y��y�K��q�-�al��'��xq��Y�&�Q����r>��(beȸ���	�ᦛ~G��g>�a|�/㷿�.��3;n��زaF�fGЙnC�X�v�����S���U<���q�ޭ�t�!s���~n�0�y���w�z>r��hN��=�+cۖ�Xq�2\|ُq��Ʊg�D?�Fێ��fA
���w!�u�\�[a }�tv/����$����J��9Ж�Bv"���e��8�V�2hG4e#'����)Բ_��$&�	��0J���(�G��o�Za�1
TS{J�$'��K��`l�S�DEM��! �
;�F(�!�P�d2C!�orrD��N��\{�G����(`hx�@?��B&�+PFa�Z٪SQ�	؆uR���1|o�8�WV��e��鞭Rk�9�*U��
�nȀf- �R�G"�{i�Q.+�Z0�:�THe��!h8�OTAU� A��V��v���.A�������g�]��X9D<; f��y�b�qh�H��C��W9a�"1��0�d�Q�MaS�Y�B��R���F�������z�"g��Ok��<s�0��l6�'q�'�g������>sv��4�W6�]���_�x+�t߫x�"zb���������1�g�V�ŵ�PYDJ�����B]���5�Z>�ӊ�(�¤#���:��-��1J�P%�9�YQ3�
qnȰ��B��3�{�5�=桻�3Gv2��!̞�š� J��
;�ĕX8>
���5s&1&�7�^�SOZ�i����kocš�*h�q�Q���ϼ���\�C۬��:҃�5���~�?>�o.�}��[�o���t�?�E�����d�����̪�_|��@�K� !(=��j-�����H�zhM���sOïq/2ͽؾ��u�]hm�`�1���?�!�	o��/���]�x�ŧ�eK�z5?% �7��G�������I�(nOG A"�ds�l����>�U�	T2�V��ǓN9���0bZ3�c��]�e|�W�g��!�/�)��?�y	.�� �ϯ��g��cU3奄�᷿�37'�Ħ����K�}����~ժ�q���ý}	�n�0��]_�����/�ŏ~w-:x1�9嫜�V,�Ӌ5�v��<;vmÃ���1ɟsW��25Gk6��_�X��D�>I��c����2A֎����\�4���L�������2�Yh�P�m!�~~ƭ��&8U~�LE������ڱ~��s]����Y�k����^,�u��HČ��ɛ��'JvǱ�tw#�F�)�oh0�R1Oe���&ǸI���k��sO?�,Vwvoی��bī�&KE�V�eat���h�~f�1g���/��cOD!Kv��H�9�(��2��@�ʔ�-*7�O�d��*'N'x�* -恌+�IMI��G� U�١�v�of������$���]6�H��ʿ���ʛ�˗c���2�Z��k	�Briu�9���+X�|�+VM�J�J���;�~QN�¼���#����3�I,��ŧ�s��'���`td'.��$l��"�ő�^[2�+���]��f�j��'���������5
�T&�HP���ki*ʚ�d]��3k���.LI�\��s@)�u�sC��ёٰ��	So� ŅU�{e-�)��!JL\k^��H��Z����s�G=�V`ۦp��e�e;��ĦM��u̝9��#K�/��_�|��N+r�a�P,[�ĥ��%8��;���q�"��λ�nB/�H�@,��`C9��G^��5��O8YA۫Xho^���]8��c1w��N,9h
�~����ޒ�{/�8$Mx�5���>�V �	�5�H�{��;;p�ҙ�h#��~sf��o��@��,b�6�c�'y� z-��i]��v�VN<M]2ĦT��w!EP}��g���aGFqϭϓ��I�Bm� &���;[Q���(&��ڔ�mD4p��~L�ivb\G{��P(S�'���?�}ã8��#�s�w�2�,�	��斯��?��w�ځկ�c�̅�.����]��⏷�
��*�u�4�O\�~���9��ų�=�B�P�P��sϝ{ �9g"P�u4.��W0�����k�t�aش�(�������?r$�9�|�����}�U�Ζ>^|{�;w1V�/���{p�񫰒���{�R�m�R���0�Ț�d�(�*ܻ�����J�`KŢ�֌PCTq�a�Re+��7W�oh��ncdhC��6s�q��G�R�����{�����@ߐ�s���|~���B1�C*J�-���M0��MI���+H%�x��ɦ����H��ɕ�%Rh�4ah� ��â%���EeS�A����w�����҃�Fn`vR����0-G]H� �\PT�����Ku�.@ .�
1�� ������: ����V�֨ &-A!IK���QFo��U�9O��՝�p����vcf=D\ ]\A�H-FpsQ#�Xd�!��ª�l�B][r�����QW����G�@�m_���[��U}#��5�U�
�ZT^� [��^�l@i���� �/��|����>8Ě�0�-y���­w>�huf͙���r�T<w�ġN�k;jQ����������É&���֦�]�Ė0nK,�7����Ԃ���¤� � �(h�ۯ�(U�%�a,\U�ưw�k�;-�/]r�)��7n$&�Ʋ���Zq���t�hJ< *��*�4��Ab���9��y�>p�m�#������1��y����{�	�p����GԏG�uce�ݸ�/�ӎ��n�BO�7',����g������N^�SW}�&37b�F�+`�@3�p�Q4�u��{��/�4I�Yh��o3
��8����Ꙧ��;�z�w4FJ��M�m�:��X1��c��#ś���w�{N�wϟ�~�	��~w>�v�NR��(�[��a�"@�d���R���g?����Y.\k�چ���Љt���OmA{�M�:jy��`}��s�ᰕ���KOB���5�{��Ep�1Q5J`��N�r�q�������7��>w?���d�.�m"_���2ҙ�M�Tsuט8.��y�G�Mb�]x��������f�)v<�f��>u�r��.�Ɵ^�o|�a��iYHpJL���MM�����8͸,�.^��+Ap�s" �h^�*�$Y�D���&�k\�H��(���!b�k���ʥ�����XT�-����T�,�D��X~�ȹ��93�:d��V�0*��	 �1�"	���^|EYW>�ǖ�[�d�Bd9V��$��OE"n�p&a&�`516����n��s�b���L%�	E#�H���mTU��ֵ$v��Ÿ!��gy��ˏp+�_�\���FS����N�-A����5B@@��%l��?ժ�s��u��}*p���D��7�-�)�/	ϩj��\��s�A��
��B0J��6C5O|Ď��Z�k�ټ��	,ȥRA���#�[�z��Z�\�8�ZHR0sgw����{z��{&1�7��g�����B\	�����x
Ď0y?�0�F+V����QÌpm	�9P��V�����fA�)�x�q��@�/�[Q����Ϩ[�Gԉ��q�$l�1/S&��'I��=g��R�W|��C�>?I�cE�^Me�l%����^�ջ@���+w֜6�A��d	�~�w`�x��G?/n����W����7y����[B۴6���p�r���Z��s��k����:Ml����[�m%���s�8�}���O�O_s2?����}��sN���`�ro�3�<-M3xa.7�C�h�`��Ww<�:�ĩ�\~�Ihm���l���i�,�}��DW.��|���׬�8����ˈףf��.bM4�� >~�m�aA{�k}��t��q�P/6�E�d������x���X�԰��}�4�ۿ�H�E�@&@�t{�L��CDIi� �6���mRAq��ҲU;p���g.?Z�n������3W�X�C9ׇ�������)Ц߹rE���d�;e��a\��S%C����cެ94��S�'��sm�2y!KY�����L'k��Y�)�����S�4�� &�f� �+�KI۳g��|mmm�t��T%�"T�V��e	,!u��t����L�#����	z��������S�6�pb�X�����t9Z
g��=ضe�F�ZB����[n�X2�l��n9F��p��cQ�J�d'��ba���(4q��	���|.o
#���و^N�t��׭)F�N�h��X�n ӫ����wĸ�%���?���︆�������`���Qf���7�����i9T]�c�%q�e<!3�*e��6%�`�ˀ�}Q�2b�t��R%,��JB|
ͱ����Qؗ}�T,;�M|�+��B2]A��+����������D7ʅ"E�A���u���Nv+:F��ٚ�"�ٮK줮�!���Z׏��ĥ#�r�b!( �R�� a��?N����7����U	�h�ޙ�$��m��/Ɵ���L3Ϟm}�bT�	�8�jEaGH��UL���=Y��U�XH����o����������0Ik����3��s�����f�I`�V�Q��d6��7�t���S��ڟ`��������FVw�uW��g~�l�Ho�/���/_��Mkv�U!��,'��Sk�_Ȭ�>�<I���o����UA[�6�ާ�{I���_>O>�k�g�ˤ˩+1l����?�$����[����7}������r��1�ƱI|��� N8�K_��'b��Q�{�[�����6���>���,n�8V��Ã9,?|��6cn+vn�up�����;�6��m��(��q��+�UlZ��'��K���~�����T�鏞��?Z_۰��_x�,"wM�
&Ѻ���B�׻��Ƨ>{%N<r1n��7^�E�:�j�����g�ބ�6Q��۷�D)
K�S�Pz>w�X~H'�8wc���5uM6uS���=��KR�ć+A�)_.YN�\%�FȖ�ܒ�Ձzlx�s��>+���"���?�<�A�����5�d<����0���NKI���d�c|����x��5�h�b�CZ$�t�A����z"e�C#)NdK��݉��� ����fl�[���Y1m�6��Z�1� 	������I&*���m�K�xHl��|�"���o������J�T�h$���~T�Uj���8�pIs�_�X�A�S8��Tn�a���[�6�=��/;Ed�Q����s�[u�쐳(oU��;F�r���}[�	�l3�-�(�C��������._�}�KW�k붧!�5��-ZI���K~B3=��6��o��!�AY�yN��l� ��
8�{&-�n���,�d8�� �@9Y^��l<�fb�lZ +����u����i�G���ƊT6H���I�T��P�tdl�$oX����� �\�Gb�J�q��K�x�,��Ǉ�r%�4-���-`�u�ƕ�a��m������x��!��g�}�|���Ȅ�7^]�E�M� -ydi.K����
����p��V�������3�L�u��y���,��/����׿w)��؁3�\�7���T/@(�O<�==�zg�����䄭�q��8� �'^��� ���#��F��ǭ������'����n�FGq<��wFp�V���}�|���{Н1����|��gpJ�����:�<��Xu�r�y��'�+8萹��g��/�{��U��1��~�m��-�8pf��_�r�����D���`��n�q�̙ǥ���~w-4����"YG��t�p�yn� `�X+N��:}�m���z���Ǧ�)����)�VND��M�"��8���a�M{�)Ѣ��+Y��Y�� ��Ę������>��U&
���sZ��eG�2�P<� $ %VG�P��/6G6_�5
	C�6��$馴�{q�����K3�,�U׀��&I��K,���TP��>�ZD�З�\�d^t��a�V��&��7l�}�,}.�L�PG�I��B+�!���~�2�dOXV8P^5M�����mR��u"i�*�J���3�ξ΍*K�|Z{Δ\�]���rX��E,�P$$��Ub����e�q� 2�[& �Y2I�Sw4��x�a\'r-��ΈQ��;�˫�8�~�j��)���Q*�眕�꠹ښmU���m�8V�o�ߊ�]��N]��^�>�󽓸���:���C��Zdغ�#W|�N��Ӥ(�5[q�Ta�ѶηG�⪕��x�K�z�f�dJ%. ք{#���Z�ѥB�H�ꎢT���-y�QG�%.�|��h�������s�QS����qkyUOs���&��u�����h�Y����"��C ��=z�|\�ɳ5S�+ӄ��1lo]�^Lf_����%�����`-��ҏ�ޙ���{���[1��94����E���;���/�J�5�I��	���x5Ue�V��nj!v�r���.I�?�`�y����E��?=�������&�J��߾F����R�o����2���ѿż���^�f��i��P�Ќ�K��<�sͼ|i��cZ&x�M�᏾��~�~����?'�s ��G5�8K�v�	���oh�ίo�"�X��)�Z��\�ˏ����h��ŧd��z	dx���#%`�SE#��Y',�#���㎞#^g|��⊫������4�bD�~�R�(L$ňETr�)`�L+YdyJI5�d̩�1��r��P(���Mo�<c�s5�TK�
v]]6���Wjv]O�w�@�WEEUM䞂�y�@P�w'*�Tt�)"��;�Ŋ�^⧶�|��	�n0C�ήv����i�� &&'���h2'	�Zl��o��]��G�|�R���UM�hkƎ�!uy�&Kd�*��<��p
ک0d�V��Uàe�$B�D�.Lvi�C�14��g�Y��0k��K}� �5hh�S�I5ԧ�����uɻޏ�r^�n�*˚bת$�D�p���}4`��G+�}5�ɼ"�K7���d!6/�LQ�/T�7�G@[���TdLS٬�C��*e���ѵ��w�@�I^R����]d,����h"wڴ�2
��x{�6Tr��C�kS���DK��G��X`���#!P�J�p=	K��ZB�lS�8��ʛf�H���\�ۡZ��Z���e��RX�����cw-O�w~U��F<I���!�&VV��V��QB&5Q�7B�V����
�3gN��!)�������(Mg܏�|�l�v����G��:z1�y��س��,'��=��[L�w��`=�-X�|Dъ�U�������|W�;��)M�a9Η�%���<�<����������4�y0v�}�wR�~���=9�A�M��/ù���߿W�"��W���6c�Lcz���ڤ�e��\Pw�I�>Y�]@��g����=|�&lٹ�@}
�:'�e��
�#��sR�͍/�s�RC{q�/�����*�����.�n��Wx��������&�l1�fyS3�&�zL��|�<�ṗ�����i�8�.l�Ϳ!������.4u���d	�14��CDl���O�!�|ɀ�E+��$������L��4_KO�/�/72o�FF������1Yl��JR�_�ŉq
����xŧ-`�'��Q{H�k*��G�9��$�����$��C���l,��(Ռ9$@�l�ߢ���F't��6� �2~I�r�)T��ꓖ�I�ww`px��_�D�(�D"��v�B�k�H�H��&�ٕA�%��KM�p� )�#���eH��T��$�D��
��o�7iS &���X@=p�́q9.�#A�d��6���܆i�l	PJf���$�B|�����\�� k����/\��~���Ca싁J0<��7�����^�J� ��G��W|�z<p�g��g�z�j܋�����a�X38�~����.;]S_{���-�4��D4�����ඤ��0.�j�(K' !¥9������K�I��~&`��9�%rEQ,i���r^M�彧���)MѺ�������ՔD��8�	���Er�(�퓸JrG�R��QR�V�VNua��8�fOt��k�l���?Y�����[S^>kvxJ��M�G��l����9�������;��[�q,9���	������Fc�������g�z���%�2���vg{�������8&����!$�R\�)p�i�WJB+K������])X������;C+%G	
F8�J;ߘ�P"�S�r��&�A:܇+����/"�9>���,�'s�a��'KH,��8o�{Z:���?{4ڍO9mmZ�qъ�\�o�׿�Ƀ�������x
]t~����E٤ĢC����|�"��\�k��,�����L��5�z��ܸ�z�R
Hu�T�\"4��bѨ��b���qD��("�<5� AY.�-����� �yD��s�	!IsjmN(И�_� E����C��݊���0�%���5���&��8�)Đ\�D�s),V|�R��~0�`�QRt��pD	��XCd�X����?W��%���GШƖ�^{�)iv�/0�;��B�5%�r����-���L\+ޢ��j��O�TsV�5oJ�兊V�I&N�.k	7�
׸Nl-h1�[Z�'k.���P��,*m�%k-y������$3(���\jhqI��D�cj���v�Ӷrz����YK����� ���U5˸M,E�ljBn�2�J�?�q�
>~��_`V��+��4�ȯ}��(zAVRb:Ƴ�GOSvHr~o��"��%�hM���5P��B\����>+E2v⮣�T�̃�)�V�;RE�sJ}�0���4���Fy͍��۟?��VG��D���ŗ-� ��T�:R���lu9�:%)��k�Tު�����4�*;"ش}�M.�L�4<������n,�Ջ��R3q�^�&x�I<��Z��b|�;7$�0{NT5U.W�C >��oa��\�����;��3���y��첕x��<v���&��)�"�`�^��V��W"˹~�5x�iK��_Wc@rm3m���� 6Y�7�T&��]P�\�����ꛑJ�8>Ii�C���l2��l�(�W���V�)<������q���C>��φx�{����?��J�hǩ3\�.����c_2�)jZ0$���yLS�^~usgepǟ�R����W���PG�2��tM�0�A���b}P���b�QP�$h�59\d�bR_��hvU�7zM�u貪T�A?){��Ӵ(��Ga,���@(���0��ֶ�Z+R��09Y��~_��,u(P5�<�&bܨd�Q3^qcL���ݢc�4C'�� 	j����&�Z8B@��,�=t��`۶]
R����	�.s��:ZӐ��XԸ::"A[G��ö�4c�c%�THaMI��|_���l�����^�#;0D��H����$DD�/�߲��f�Y&��l�z�z'�����JNs}J1yAП��?�9�� p�w��N������Me�h�o�ѩ��ƃ�k��(x��	dK�\�� \@���N�0T���G�Ț� /J�V�U>�g+�Q*�h�T��{��G>x�~�k_�>~�7���~���ࡇ�v�wY[~\�{���*Rm��K���8�sY�le�5I���E��Uez�4�]�Q]FZ� �P6�)0�ؙ4�A#��������>jk��l�9$�댢o����a�Hd�Maʱc�*Ѿ�Y��!�1͚#�-]GjJ��=_ʔϺӂ�^٤�eI���I���'_�s��i����l@��$f0w\�2���sp�����t��:6gf �q����ﵛ�(`?��[8����wo��/�h%n��TYz�v"S�Ѽ�V\\��=�9��� fϛ���3�OC�?���?��{(���uz9tO�ƃ��F�y��k�lܴ�f��UhN�#�pLG�%�A��Z���om���n|���q�r��e�ٸA^�ߍ?{B�M'FJ�p�oB�X"��㷿~��
��7/������@gO3�ۻp��AK�����R�ҽ���=�i�N}���_��/X���Q�]���9w��"��ID�	�,�Hq�rpuq�(0��5�*U��|���|	��c�,b$S�""�!��t:izK�lmrS�@���8��-��{$�CR���i�t���Z�i&�O#�Ik�z|dBSv�.+�"	��Z�'?|��o�駯T��ʺ�3��g�7M+ KE ה/���ю];�`�̹bP�4�%��Df��ӆ]�FU��5��[�V�h�$|�u�pS&�tS9�"�6�U�j����D�TJKՔ;K{Th���f������.�1d�����ߨ���+��W��T�Z`o�~2X���N���#0y���G	�ma�Ņ �۸F�p����e���0H�5������C��
k	�
�Ȼ�������x_ykGq�����/���q�+_�f̰h���G�~��pӯ��zva뮭 ��N:d�MJx��Қ]V�l�$��Բ�O�� v��ֵw�}�$�'��r}ϸ����ȹJGԐ��Ѭ�wF&���&vp�n�C2=���t�J�}K���~+U��|��%�@]�y;VLMrO+Z�sĸ�h�v�����4S̝��#̋ٴ�0ᱱ?��L�/;���;��9����%he� ������ �7[(�nE�)Jf��������k��Z����|����Y��� �M�x�$�M���&�v�~F�������1��d%U%�I�G/�����v6����w��7=���Q�趖6�b]�PU#�a5u���Ƒ���t���l����F�<�VM�-�L���g��+��ݷ?�g�݈�O^��ݬ�G�p��o��1�q�c8�'�����ǚ�T�����ʫ���Ø�3۷��/$#��'��rn7��	�~�#8e�Qڹ�'��:`���Q�b)P�xV��IMU�A��xM�2�DHz��,-�TE
�LpI�^@�T��J�2��N��>���Q9U	`t�V-�g{ʬ$$`5<4�]�wN��Ș�M��9�W}�������L�+B��4=��P&菌�{��Q�}�ITZT���,/YǞ#����h$���A�"�C**mkCjJ%0�G�ój͈��	��<Ʋ��Z��P.��!�]*�M��ي:�7�2/iU�La	g�jyү��oԻ�*A�A��l�}�fɏ��|��	��������/O��߽<g\1��.�sK]�(X`���������!�LI)��!a��*�
�4�`T�M�헻�}Gr:;�y%E?6C\��>������
�=g���?f���h�M�աUT�fX-�p4;RC�$-+�3/Ʋ�t���ժZ�ڰNj��n\����բ��F0�ҔX)����JH�ô�&�qt�jذ}瞶�y*'ZjMn�Ą�j	j8�Ć��� 
���o��
c�T dK��F*�C�ĳ94	���Ȉڣ.zz�R��a����Ib��1�ܥolmk'pN�h��_-�,p��^*��Vn���J ���Yu�&��F(YVg�����XĘ��B ]k�i��h�Hj[�^�_+!- +W�l��f�d>���y�^��d�,I���6��ؚ$]؄Mi���+q�zP���m��_������%��v�_>�����i.�)'�q�u�R�K4�\2�"��q�[|o²���q��O`z�|Z��=�ݳ��oQ��|T�s��p��G�|����		���y��	��!qi455� �KeLid$W/�i�Ĥ��H��s -I.{Ӱ<��Dn<O���&��hNA��5M@L ?i@MK{�~�v��'l�F�����3���ϡ�df���r؄���:�1��ͼ��Q<���ɤK�</��H�V���)�넱s�a�¢���(E@r�߰����l�<���X~�r,�?��V���[H�������xȀkA����;��[obڬi8`�<m�Ow\<N�^�'��f��q���84�W��BT�e >�r*����`���cnT;�����8��FBAբ�'r �'B^���� kY;\V𼩞&�o$/[����+F ۤ/wI�����\e[:4r�MN�j�����2mX0{6���S�4��ҢCqk8jy��$X@�w�-�`hl;e��:�atl�rg�1�N���*.�'(@�M�YpH����@���(i�%J�v�f�Q,�DL��D�����Bv�Bs��$+f���Jq���BD��E���"�i�?�^I���o�NFz�<9RlD�)��ؾs�>�����$�dq"b��V$��4�&�#�	�R��:yG�x�+���	���H��O�WP�i�O���ֶL�Yn"g��H~.��r-�6�Z���}�ʐ�tP6Lm*ޡFNp!e�KE���2�&}o$b�"����kr� ���,�|�*�$���5Ⱦ׉G OPy����Q�%�ESwN�l�]B4,�͠�ī�D���r��#%�==3�w;s�\��db<�Y�(�v��0���7�{�,�M�0h	�^uc��EE6�0ki�Y�֔yk���lb;�J�7g�E�����ako��T�[���%m�䖎��iǻhT*�l5G�g��M
,þBa�h;wД�����={q�g�r�M��J�"���2�r�yrʏ����q��!��YlܼI]�׭��Rޢ�I*hwwwb���������&�]��Ҝ���K�,��{`N����$�+�>�*O�dZ2-ػ�O�z�v�l�֣��%�P��Ȳ�b��H]���?6ni �V@0^	[n��U�?�m�����_k �?:�%c��7��G*Y�4x�X�ȅ��ĕf��l�S9�њ(|1�	b�7�ʵ)_���P�>�Z{n�� J��hu�:����m
���k8�C�b����Y�ؾu��Kʫ��$#���۸��V�������{uZL��(�g-x&�g��(D�������T�`[�7�^#i܎N�SV�~�Ȼ�i\��Y)��e�~�0�/��y3Z!�T����JνW)���܍��`�T�I���T>�!O��(�_cm�S7�}d-� �h��+˅���\��*�b���aR��im!�.�hNP���h�P��x�-� �k�kdqBk"�4����)2���d�J���� ��lJ�-CS�+j�%J�~43���$���X8���h�*�p��T5� 4�8�� �F�����E�	 �9CF˅I�k��\iiI�����8��v^K��� H��8�f�P��B<��t��"�n�r�!�""�[(a��Rkg;��M?�#є�xQn�����E��8�U$y_��mش�W�jX��L*0���4km�6����1lݽ3��102�B�g�F�8t)�m-�.(��I�_.W����Ȏ�ע��Z��6�T
�L���G1��C�*-�-��DZ�4��m�߰IKͷ��q��Mvww�9c{��I����9�lvR����H�����w� �@�M5�e䜆$�?�q���c���@i\�4�Ջ�CkK+bMM�6���<Gs�KE�e�2W�_�?���%�[Ƅ,M:���q��b�}�џ �gR�g���qy�n�گDR�����ZAn�����^���K5,Y�}���
�˥Ͻ|��8����3ےV��*��ߎ4���$uԆP)�O��l�T�es��W¢�3p��#�Y��)�����{e����O��������٩GL3�����sZ��8�<�� @򿤶=5Gz� �m�\��]�
Ka�L�rj�W���w����"�zm�|��7q�U'�����-����B�ſ�ؾv@�,ʬ����k�r�/IRЩ���~��܀�~m��N2s����Z�j�,�v�L2� P�5rF���0�GX��s��&Q�J��]�&O!_�d�����:�&($ѧi	�M�&�&'G5��u�3��eU��D�\S>��3�wUD�i�A@Q��~`�f���7�O��Ԇ�5|����|��)r���=M��
�Ta�d�b)*��$��{���;U�ue����:���V���x��΄�2�2��68�jʛJ$ni�F1A\��h�GS�p&�&Ū	�y5_}�b�U�
49�0"?`E�eX��D�������{J�e�eSs��H��#i�r�AQҳ���K���SO8F�&�ʑ�;�4E�
�6��k�t%��p���xy��&�9�Ӻ�i����2�#�`�Lf�
܍���;�z1*��.8 ��*CE��-?�ޘ�h��"�ʝN��陦�i����h��o����Oػk�;;��XF	ڔ4*&)Y�l�~,X��|��<�x4�e�:�׉K:�t�p	��v�����Fsg�oc��ް;�	 #d�,���}.�Ft&�5U��؍���R�d���>��_�@�En|�.p�J��b��n**C!��QE><gC��zㅪs���Չiz�h9�t��n���eS1���ql�)܆o~�L��#�\�C��|g����k/n��H
{hmi�Ȏ.�m�B�X�Ĥ
����Qo8k�%�Q�zwm1�r�)�+�+�Q�}�o�iF�(%�����KC���^#摪���7��h�q��ñ+fb�¹p���q�#O�4"7[Г7�UY�a�?D�&P����u�^�UDiN�$H/�:��]�B)���k2>mISi��m�5����T�o,���"�y%A+�{Q)l(�(���+��~���M��%�Ě�/a��]�u�g�q�Q��a&h��:�%�z��M��N��#O��e�� cH�ܰa�W������&6�dH��5Bo7�ڦ����T�<Z���iɪ����7�Ta�W�=S��7͜4ǌ�w��!^#.M�0)�c��8/��ǟ]�>�X�4����8�^��K�R��o/&�8ҤS�?�1֨u�~	jב�ǔ�I���A2pT�}Eŕ/������[ūj�q����[*���9ӻ�~�f*�.�I����ө|�Z�(�<;�#PF�@F��:�3G�I�Z	Ӣp]s���vbV�lDSFG�zM���.K�Y� ��gܟx�A��rs�1��vk���q��d'��~`�q����[W��Y�����ػw7v���'����0:{�c,���wl<o�)$p�G���=`���9H�(���J����\��M״��q���q�HF����z i�$�k�������}Ջ��Q�
m������i�����~���Rh(G�oO�q�k�/�q�T�3�Q��i2�>ր�nL��|�EX����P�CE�JUa���$�to�3�ܻKZ�{�0Q�_x��q*N�e8����3r��hM4�%˩B5!��ݸQ��Z�v0.Kol`��2�y�Q�\^׀�Xz���I��Q��I��TRL]�rH9�S�˥ZD�s���;�5lX?�-����#�5Y�$>-o!�!ӡʌ�nk ����&!����ѡ��b$�c$QQ��1�������uSdI2N�h����ǻlp1��BG�*�*S"ݺr�	�,Ǵ�8�4.|סظ;���!���m���'/>���w��&��� �K[�a�0�B/7��A��D��~�e�k�Vj�c�t²�MHP@���F�al�Jd��g6��`ڮ��J�[#Q��&	�rǕ�I���`&X)����|~�nr7�u������]���$ˡ��A�<���;�2��̙��5s^{k����(���ķ�׷���LUaI	rLPK�3�\�מi����Z	:�Y�47��]*���EtZ��NK�D�J���SR��֐��&��R	���$��C�bF&���9��ao� 8`��c�I�hT�V
�ܠ/C�kT��CWG���1ĒatO��JJ-�)���,�}�|�̭%.#�}
�a*�SN9�ϕ��ю��ш����B��~a��ȿ��U���C�6�W����V�[�e�	����Ұ�& �Y�H[��\�O���+ڜ>�j"[�hJ�B��.M��`�g*C���W7)��0v��Z+�y��~,֚����Ӿ�%v�3�qY���v
�W/�u�0�)�2�t���`���Ov�wٳ�N;��	�\�R�(�ǍB"�_�D5f#���v��C�EȽ/��<Q�m^�kW���&��G?zn��v,Zt�}e� ����8��לDM}ޔ"�?��8LV�A[�٪��&	u��3F��Ae�)�r��a�)+�Vz�Hi� �X�q��%6����w_s��9Gb�*���I�� k&V�K�\0WNrg6i�74���㏽cֆ����{�:�2W��ͷԗ�F�h�Ŀi�L7A�L�-&;kƬ��Fp�&q��F�?f���?Q;�d�Ás�յ���a��z���vݖ1����	�>�x_��	�U}�$��fR������՛t��������i���q�ܠS\���� %YoQf!f>�'��'�mt�Dx�i���X�d'�~<��8��y�1���~�+p������Zy�I[=�&SN	G��-,�R6�	M�){�i�ų/=��x-4�y�,X� �AQ])��.o���g�Ծ�pa>W˸�򥪦3��g�CF�xTRqn�dܒ�'�l<��[JI�HaK#�c�Ae�m��6�Y2]� :n[�)ّ;�U��H:���"#��5�T����w�d�8W5�_767*%Y��J.������7DI%R��Hq��T[{�;Lzd�%RRא�k��ۉ�XE7�����N�U!H���W�]:
PK)������H�!��q��I�`{�tif��O]�=�7���-�D��k��(�9��S���2ys+�	�r��a��}թ�A�4�Q���T^+��������o}����2M.���/^����E�B��;3��Y�1w�t�	FK{e���r�|�.<��F���%�"j��>k}�?���>7>�[*���Bʭ���I���u۸���Rd���xrC��"�LG�n%�����_���zu��i��pN��o�e�f��i�Mwi���+cص'Orԏ�!3w�^�)ֱ����0Q
e�m�]9H���I�������e2�P}��G��#8h������4�L�ڝ.#/��pU#˖�E��]�����z�(	bJ6�}U[��c`L
H�䖸i�PF����جr�T�QU&f�4@�M��)K2�w�ҩDX������϶�Y���]��w�Xr�\j��f5���C>�����������ݦ_
�G�6=]i�\q z�=���0Y��e�ҋ#�i3e޾ɋ��PP�936a���A�nk@�`���=o��cm�T.O�w���FM]a��K	���I��
7���P�X7=!�F�m���#�M�hA����9��#ҿ�ѷ��N�=&��Ӟ�n���gS�U٘4ڑ��TSʧ�T�Koa���^)5_>��=��l�)��%��\PFƲZ}iU��tJ����>Y0w�iN��2���&740�w<5�z���c*��;M�(eݘ�n�4H�7�+�)���ϵ��5pt���B��T)�&Ŭ1_zI�\�)e��/B4�"��~�u��U��,�w�4N�v��?�N1њY�FkyN�,�h4ETuh����ʹ�����
�Fш0POzv��ȽZ=ss�I#�߽�v�}W+3��'>�n���O��N>\]%%n��]�=l�	�Y��k�G"��rY:�����A��$Ι�ˍ���
�tX(^mm뙔Lu���,�(7R�A����4�$.����*r�qZ�E�	�w�Bss��%�:v	n�m''�#�p�i3���z`Vo؍��?�xX��r�%����o"hͤ�k�C���)���{DLsa�b���+m2U��s��7�DZȚ�[������YF��ӌraLߗ������y��1�����O'C���ǉ�&�uc�I��A�����ѣ�>ֶo*蠦�y�0#GM���������ʫ�=!�-M��i	�Xv���Ԍ5�������Җ���V��!�f�	��-�ڥT���x����=h	�{��խ�{y��m�=��T*���Fb��
d��ʬ�.��,��^9�T&J�EOw/6n݄M���	��mp]ⓓ`��a]�u�
8�*'��mݷq��9 4Qr_��z�YǸ���Ѥ3_Er��rK���&ƌ{�����GU��5ӑN����N������:���f���y)K)o�eԦ��(l(�E�Qu���]��Ay�%�(�b�\��r�m �Q��F);����x��[$�е��!�|o��\��m4�w�״�j���I��ȒK�!ma�|�f�8!����3�F�e%)~_/�:�Tc�)0`�VP���߀������7�-d֣e�F���d�ԧ"���kV3	�SQ� 8ڰ6����Fj`�����';&k)D �V���V�1W*�1{�A��-wa��V��?w��x��8`�LM-=��-ذظ�e�[f";1�dS�ޏS��	��U������\�փ1AZ�ص�іֲ�@ތ�Qo��n�ֹ֣\��db�=����3�:�XR]?� ��/pl��a����;��H��avO+^|e3��
_KM�v�,[ڋ[�|�.��w6k�C��k$#��^�Me���n"TUsO���I�6E��풤?Ӿ����a��I5!W��ͮ��V��<�R%�c��_}���5Y�-ӌ�4��"d�|�H���!�^�-�fıf�)�2U�	�$�7�����4��T?���qE�+�_Д�)�(]�B�L�n��	pHɭ�&:ξf=�8ѭ����Ncp���Hb�u�|ar��3�8��Sv�t�e��ڂw�L�G2�F��;7�#�M��J�&%�r�A�A�s���iJ�y��Y���:i�?h�B�t���uU���ߗ)#�	W���z0�ҫ:t�p󽕫:Tu���9'͌�H�%!��A����,xXF�	c�`c�0Bl?��B��@a49OO���]9���9���nUK��5Ӫ�u�9����^��_�ھH��G��#r s���4Z��X��� ��v�B����������<�����Y4�Ѭ�+0�i��D/����N�W�������82P�f��o�Ap�&��B5�Qϱ ��'Bc�#�$O z0�G�l�FF�A�,[!��l��3I�U,�ĩ���Xz�w���2�;�(2B-S�鱱k[.c�)6��ġJ�3�c��w���7�H�[\9�E�A�}��vRw�1�mxj�
0N�#�.H��vb�&l"��ԣ$��?9��XI78��%�����y���`N�n��������cO=&O}��#s���daiM>�џd��n�����sյ_�������i��֍��b����{�o�ٌ�w��V#��T.e�h�[n����Bl|�5��%�@M��F:�W<Y���H[4��l�L��)9�R?�?��X��:���dx4���bF%O�:V�'��S!���|)�{�y:�0�K�|X�P�<�����k�29Q�ne�y�ȃ`��V7g%� �g7~���r��l.�>�={F�n��:�>wVZM�==������7d��Lˁ��՚����"��$r���řQ�O��&�2����Mp���@
�݇�Hmz��Xc���A�n��
9~tB3���*hvb���'km���5V�V�$�n�f�*�������CQ�C&��_��{m g�XAS��t��<M5�A&aJ�L��4&&4ż:�PHIG��댌"_*�l�L��z�I�`��H�Ux.
K8BM���F�y���F��wJy�桂�2A�CU��c8��T�5�L��"���A�F�;�5M2��M�M�F������*e���\�4
rι�d3�0���bK�P���æz±�Y[�俷�V����7�u���hT�4�.��S��|B���\,�NW.�еר��Q���juɍ�I@5r߸z#����p&n��x��4�r��=!�׉��v���\�α�@3���K!;%�˚l�F�чɤ̽R�}�H�zV��]a��Y-y�9T#�#�Jsp�(�'H�ޢ�4p�ek����g��N�7u�[2V��jN�^��=.��{��\ȑ+Y�Q5ب�,#�HJ)��/ȯ�������_�(0�7hgZ�?�g�(?1�\L�b<�����IObP���^�T�n���T��$u�>����@R�f��b+_��G�WoWe�`�V!���ΏIO+���Y{�Q5��X�mo�hπ{�l�H18W�rP���C�M��u����X�/6|���.2��to@lw�h^���-n��4%Xb�P�nAM��M�~�}�I���	Mg5�=t�"y��������1��6:U���$��zD.̓�$Ͽ0-�$�޺�:c��MqRK/��ڧF��4o��1k���/;�I�D���i+�]H����M��4���hH��҈�j�%Mǋ�&3v�5�(U
2:���:�O<wB��x�=:)��~[��.���R,���5��ZM����R������i�+�5Z�T'7&�r��D^/�S.�H���j]�z�:̈,}eG�{�X+'n�Yz܎h�a;R/n��=�Z�)nlե8XO�Qi��~
�[���YYn���D�nޞ:D��hzΫ���zt�c�5���V=�Om�e�7�'�Dx���rG�r`�̀Z��Gsr�ޢ	����zݛ�[���~����^�o��H'���"çNϲ$B2��Հ����$'_{]y'�����+if��!?p�E�1
�x�қ�(��M�-e��A_dC3����xx����y�Q�7N?�PƉ����{�3�n�D�����2��C]ì��H� ��)N�Ov�l�>�a/�����Z����3N���N��{U�S�ef�￐�f�ْ�p����w��g���?ɧը�}�����|�g��L�^LޱKH0�c@o*6�i�����}M���d�)֚|*���e�`���6�7��p>���9a�̦]��J)�2/H�Ƚ� 	%7P@�jd��O�]�K��lr�iC�@X�˘�v\N����j��lB!r�Jb�1c��kt�~b�(&�(B�01�1�
K��*�n�7?d� 傦�9]Sl��z�ua@����A"y�N�|B���w��Ȩ�g[N�9/Ǯ8ʩK\��>#�Ϟ��o�]�cWk��k���SϜS���6�N�t��b����0]A�)q�c14\���4��2n/w�H+4�s���n�|=p1a`��9���;d`�r��a� ?l�w���)��M�_���.�����[\���S�͌�kFӚ�1kC=����9��ԙl�%k��dZ�Xa�p�)$H����5��7}��l�@��]�1��I�;�]7��m8��4�Ȗ2a?kB���K<\�K+z��u�*ҩ�y�J9��k~&6�l/S��-�rU9y�u9�vb�>��X#>�\� ^�j�"W;���QvԸV���h���r�u��l�Yۄ��s>k��l�_���Y	�9:��q�h6�bph������55D���CI/j�!��_��KӚ���W��[n���s�S�$}>�ή曟�$H?�K��lZJ��bG�[�h|om��3�����u��]�/ү���j:�����V��ђ�4�1��.�d\	���#&l�O]lQ�E��e�<ҿG3�q��)�`$Gd�j��yi�C��;&����侷|�,,/���������W�}�������X���3&_�ʣ2w�#��+e{M�;��]�hb����!�=5Sε�^�Q��D
�f��|o�%�`A"�d}B�4l1`�2�N��`�>���G&&GC�}��"�+O�/�s��7Y�j�s7�N+[v%��\#�^��D���y�����F��5�y>��M�]�ۦ��Фc:u�� �5ۚjZ'���|�;nV�,d���M�U4åK3]�H�V�`J$��-O<�;v�������g��3��АE����t��ݸG�׶䙗g��A�]@gS7�F��a�q��2bͭ����ٯ�5����|�'tK2ֈ��sR#'�?��K�wޮ�l C>q���I����㪇���<�蓼�/�.KKr���qS^�\\��9��g���evy���n�M�Ã�ժ�����?D��'�z	5>�PÏ�#~�d�z��&q��4,Dɸ&@$��BZ���I~Z����������[c����隞9}��h7H�Z*3D����)���kP�+b���@����������Y�;��L^u��w���B뱡�^�~g+�Q���l�k��l�s�/0�43#G��33Ò�цϋOR
~D���]�B�(�N�ןxA��nٳR�F�emm��0�Q�?׿��,�?�O���ͭ�f�!9~����J�nJ�ڈ�8�kȏ�b&�%7�F9P�Z{'Y�a�������G>�b�����Ķz��pNjM�NL��F4�� c��`��)�s/�Sc��p���p��v���N��e��&)C��k�ے�Yџ�^�Q��n�X��K+�?�y�+�r䪂��pZ���}`�L�7�_��!�O�^��`�u�Z�u**�p����^`�8�����iFU�U���X�]��:1��\Ʉ���6$#p��D�1�0�h.�����Lz2B��7QE�A"�N����r.�c��W�^�=�ՠ�N�8��({�Q�����L�g�~�
Gqh��F���q���$"PB����S�g�i��>��>�����6d�ꭼ�$M�S���Ph^���Wʫ��֏�Μ9%���(������]����< �kKRA]QO�?B�*ߌ�9�V��nk�:4�ީ�EE��U�~L
��u�E(�F¤!�!�a�ȳK)�7r0��o9Jl���3�,�5us�>��5h��B�M5%��^<q��ߕ�9��O��m]��>�z�����F�#r��7��؀$�۲��	B���`~iM���g�ٴ@�2~�l�V_���L�@�3:A���e'�c�P!�C�υ��${D�Na�	YJ��}�F�*SSS2��h��,vӭ7ə���o��h[	F�7T]�^�&��x=��xR�2y�f�?2)N���S��Es�m�W34(��}����SO>&���E\����%7\�Fj4��=�&�N�7W�Wݔ#ʅK��xOK�2��45��K���F	�\�h���9��:,���P-;����-wީ�Ā:�<* �(�ԫ]3�}SiV֢ݨ_�N��8R��y�i�xG���AI�>�8�c�8p�gW�}!	G�=+��!)��WL�	ߘ���!p��r�h2���h��Q�~-��?CTN싟REx�!����d���̎�]M�����
dI�8"f.�{��ARD~��H��G�C������%�H2,�eK��ke�N�[�f�˩F�	3\���H׿��}����J�%C�P�uG���D�ݬn��Ճ�MhDb���4�Cr�c�H+��aς2���k�l@<����-��Cr��dsxk�v�A�I j�O��>���uem�#�X���FYۮˀ�A����kH��T䎛��K��o�g�5�ז����˳A��Y&�cd�8(VW����]Po�O�>!''5��!�f��x95���|A��cLc��j����Kj�z�Ɇ���4]M
�2�@��& {Oʣ��˚�R�n��)�}�S��2�E��OW8ل .@�K�i{�#�+[rhjXf5-;|�KY (�^��F#��#4ڳ˛2T��V3����-9ɢFsW]��-��Ȟ5Г�	2���}}V�]�����0Չڻ��z}�RI�˾���l����V�D���J`��]��nJ�Oi<3
��^�G�T���VL#��'�2^m4�4"���y����Qr�6V�q�����BY�4���ࡻd������sr�}o$�/�c�c���j8JBظh^�;wZ�`fFѳ��#�w��յ��JY�6؄.#먔��,�����Ld���!x��A�ߌ�e%�f�|�x���<8�Ne]���Ia`���RƆ�C�ʎZ�&����Ad)l�*�(yd�ryt,��������<|Ֆ����ؓ>2*ve1��xW6!�h9�tRvb�E�K�='��4��ډ����nH_z8iI�;2�^T5z��+T$	�9�@*#��.�����J,��S!|R�L�����'�'�}ϯ�%T�*}�T�%�nXf���m��KA3u
��qk�^M@\7�ucsE:��?r�>��_|Yܩ��󯟗��M2+3�ag��AA{�I����P�,�Ą�#)�r�i�k&J���mS��1��Rܚ̃��!&iC���	�l&��ٱ�W���^hY>|'�\��� !{�����,!�1��j��a����oyH����AӔ�+���z*L��76���bQ6�]�m=0�Z�g��O=C��9�YX�H����`�N^o���fSn��y��
�i��H\Sk��v˚��UEK*�:m��l���Lsg7.�RQ�FY���M�(4�ߋa��U\�au"e��M������̀���_ш�x^���쮁�����%W^}�L9 3��r�w��3g�������ٳO�o�&�N���(�gԐLy�Dm6Q��<�q�m�Ҙ"�F��cT�#�&qmǅlx`�(f6֬��r!���EϑX%͖L�Ý_X�{�
��:��}㲼��G��"~����<'��i��V��3��h�>-{&KL�z�!��#�^GD��nsc]JF3��Ç��w��Ʌ�䦛o%�7z����w@�	!��ݳ���׶d��Ey��ձ=,iLM�!)���&����r�M7k�sR��R���͉�Q �t�N;���Z�=�f'�z�k���v��b��l��]VywS�������o0�q���HwT#e�"�ɘ�6�3�(W[E� ��P��WO�-7]G�	kf�#o>�!�A,�a �l8��%6R9ɪckuM�R�fM�����rۭG홋A��xꂼ��#�0P�E��S��p_�yI��]6W�����D)r�Md)�-G���^��W�����z_M����\�����ï�//��/��sE5����7��|�k��i��+G��sg�-9�GMr	wLR,S����2�5x�O"�2�&0�(-���#�RH��3����:
�H���l�@I�A��@w~Iv.,jġ�³��V�&����n97=#��F��I��8�1��> 5 zxF�1y��gl�놇�>7;#g]���쩬�����ʣ��A��޽�W<81 ����Nɾ�#�}~����)y%FGj8?����k	#�nl��k��$d��ج���i�P��Ŏ����`�>N��xQ]z�<Da_��}ddX�i�|���3�=�::M�òw�>�ԛ9rX#t����p�S�]��^�W���4�<���5�ҀMlu4�ۢ�3e�N5E���0�R��6�S�6;�p�����
5(ʘ�Օ5�(�R����߿Wffg�F&��Q�c�`��/�k�2�����iuJy���FH������zmMa=B�:D��ZbskS����{���7��{����(i
:�@����96� �F'dk�QK���0EZw^Z�Sc>)Kꀶ��= �(�~�	>�5I�pO�����0��E�>���fe�������#�Ⱦ�s��E����.ݳ��]PAWӖ���+z6��1�ճ�K���� ��泍�w�<�A��e�`����u~��,,-ˡ��4{��6��k��ez�=���)�6��Ug B��j6Q{�������*f�&z�C!�q��]GM��;�W~��?B�췼��z="�k�f.=.�+3�ʑ+o�Ɩ��M9���^K�7I���x +��*Gݼ�[�_����/I�iH>�}o�=��_�⪼���O��tr�T�6*���fzA�a�����ZBVN{~��B�l%�$1%��F�u� �Ğy�e���Ɉg	xvrHx~�0�'A�'4�H� O�#�Q{��鼑]h��~a}S�^lȱC#�������qA�������K@f�Z"^��ll�eZ���`�#��0C"ߑ��8"ϟ<)�����*�~S�Z�<�����W�:#sK[���W���WC���3��i��I��.҈����yN����(�����^��`W��j9vň\�>S$OZR���{����-KK��_w�1���YVֶ���2����Zݬ�!4a�������BvXO�.�;sQ�8<�M�,5-����2M�aU���h��J0�T���l0�o��m��Kq�~d���@?���p]͠K$Q�E��(�N�UǱ-�JQn��
 ����$�,;i(�C��jӌ�� /7�ʇ��oo�d�FH�i��Co�(�YM�nF Pϊl/8�L`e��|��dqeA�]u��L���U(!!S�*��w��x�E��eܻO�''x}�R�<:�W3�}�1�,�<�o/����@��v�SM�t���rכU����d��I@�3���#NL���y���߅����ލs�m�17�bL3�	>�\4�<'��B��iG�x}��Wx��G��z�@�f#��'�xFn��F���0 B0לf�-"+��` ŏ�ps�V
��u�&1�F���]O�Q����`$<t�`�?�����O�]�IѾ�o�������(<����sr�lI�g.JA3����F�U6z� �
��Ik�����r�-G�ŗg��z@���//�Ǐ�QF�R��w�cL>�7� 2B��)�5 �ݐ�X&�����6"�a��k"Bv��,�&m�X��6��_YAyE7z�zb�	���g�l�D#�D���bc3'�Cm5��`��֜u`5
MMk���P�_��Vq��S�t�)��z\Sc>v�U����>�r�K�����Eb��Jʓ�4����Q�ꙒLNSX_�yeF����eK=^�N�0����.����X�Q�6�r��~���ǩ"":��|(w���9��(?T)�Pov]C�x)N��������]��^�M7ex�1�M���y��r��g_Y\Oư�i�ex�F���~Y�����K|���V�X�B@�\�w{'�|J!�>�+t��Aqjl5/5��>Q�=�2��4�-CO�nP�;B��[*[�( h�Ս-}v=��R.bPѦ���:p\�[+rӝo�JF0�P5� ����GL���3�u���?y�ڌ�������i�Sr#!�#��F��PJp_�=%-ht�U��]�D��M��:kj_D��|����dh����Q�8
�ȷ�q|�!�0�c�?�M�$�U��A�􍳫�c������9`L��� ���?��S��@���~�$"�_���cZ��w�}����/���7aB��6Č�Ll���s|[V�5+��[	�;����U�Q_QQ��6�.a�G�g{荷ʓO>%�~�Y���XX�����|�����G���I���׀pQ��ͺt���!�����3�����fB"W����;*Ͻp^>�����R%������Ɩ:��A=k�4`��͍yBRW�V��ۯ��͆�|rN��D#%TüK\��A>�Ȝև�H�vM��s�^_�'��nX���Oںg'��+�?c	�$_>� �S�֢�&ʺ(-�D�F6D���ה�̘f-)UrRk��$r��</�-�Țb�ס�k��tp$�@3/j�R��{Z���K_{���*!9���!C)D_�M~��+���&�=+�5�l]A�i�������6�w�pM�1n�$_%3�ﰱ؟��u�1=?/�^3��eM�IV���%t�[�Vmi�۔�rA�]`2i�g.�n��Ƞ�̭�i���F-M��2���n��ￛ���J��io�HY����<� �O���|�p�jx�qGlӐj3���cٮmKE�)$@�
�5I��{����] 5�nn������BKkS��߮ՙ��ۍ:/^y5� kBc)RC���z�����t���6�X4����G�2xHڞM��ZY�� i���A������Z=O� 8�lD<~�� ��V�IF>�ǎ=��%��<��"��qO�&��`[�9��J+6�u@���@w� bB�:Q3P(fX>�y aᎴ[Xg� ���q �fEn�� �ˡo�^)7Gj�w�$�g}����]�%4Tm$D20�/��̔)M�_q^�ul*��"��)\�]@�w���:�$�apñvWS�v��:�U�)�Z�b�^�DO�w������k��n��\�j4W9��vuIΟ_Rý����ȏ˷}۴fv���=���w��ny�������m�q��u9vZ�L�t�O݇�%���i��_�Y��'?%���G���ܦ�{ivN.Ξ�}<�߽B���'^yE��i�
s�����F~��N�{�}�,�κf���j$R�<��:��g.��ZF;t�i��M�I?i�C�/���?2@8���
���- Ԛ�
�o�B�}�=�n�'/ ���k��$4H�=� 7ی75��C�mK�8�O�>#7�xH�զL�P��G��P�UdXX\��s��;꟯�<�)V^�'45P�BNib�Wd��~�����TlK^%�׈�%���ʩ��Z���.���AǦf��1�62��c`|��4o��|v`1��M�d	S����;ujE��Ɇb�;��pW�-��:�H��3�d3��9:���N�-8a�ƿ�(����!g�\�ώ_q��bu]7�+/əgdy�>�֨�h�??M­���>5z���� ���%M	������g����N��H�JՀ����T�G��ٜB6%}u��1�9V��+�(��h���s;�,��Zj����&W!_���C
�lǢd@��g�5b�<_�t%��{0��I�v��'F����4v��i6���4~��c����E��?�9��L<VA4]o���E�V׍�0j�������I3�=f$>��C$�_��2lD�(=��o�L�ť%��5�v2BR�����F�t�B���)��TwĦʑ�#�F���OZEU&�G@�Ԥ����Y�B�2������(~�3�O�u٣�L�� ]Q����v����a����s!i�ƆeuӮM������v���x��i9|,���9L�~�/�r��%�5{#����{n�2��1��<l�9��^*�M:Ch�/|��˟��/�(�lRTG��縷��͗Ji��}��&�g���(���r��%�;șKY.t��8س����hjQ)l?2хX�O�|�V�,8���m��2�`����bs}U�=�y�34%�36,G�YS�٬�b��Q��A`���f΅�S��bnC�Ֆ<��Kr�W���Ȉ&"�q�2 ���j��ɳ��酾d���P��iIK�c{��:zX�����>h��s�˲w�~4�Vp -�9<��Sv,�I>�I�r�i5z$RJ�Ͳ��{����*jX@����P�ŁP��dbϐ��]���t����t�ų�Ԁ�!wF��Ƥ��s�і���l���Fc[~���M~�~D+y'��9���kʲ~F�_;i2AnT���q���*h�no�uSy�G����J�ըp����4��{�@�6j�֩�?(����X��8�<C*�$��9������u�����=�o>�A�(c��EN�/)�$e�k]Oi&v54�:AΖ�ɜs8Z5T}FC���L���<���#�02|�7��9Nh�b#�V:sYN	�9�����`\ B)si��]�j�xф�N�3�{F�ۛ�*������[i!}6�(L�gf�wYmZ�#���QC�Y?oP�KY�op�l:�c��C͌�j3�|�c�MD�'�=ds��qG�*H�=8j�#4`�4bo��P�e}��}�X�Mc��QA���3qd�j/*�b� @�?��?�����!i������x-K�}�_�3X��}7�ِ�{��������zϷ��|��h�
�I��.9���7xV������j)��΋������]e�DPA�(�G�F0�+���3/�K���m�������!�)�3���ĦNS�qr��ۥݣ�I�5"�Q�m��Ⱦ
�����2�.�j&d���lKeX�[��0pE~nA�f;��j�� (�/Ӄ��v^7.�Xl�A�*�m��5����ܮ���Z��H5�NU:�鳮�������
��Q8/�^�({db��XЭKe�=k��n'z��[k�-���ss2;��
�r,v��8(�w�E����E䔤K��4ºF���7%'�1���}ff�n�	囼��k�pQ���~���VCf��#_ɱ�����h޹��%/<����mo����]y����k��Y�����~gK���T��(��z`)d���T'ЕiM'k:	c����,`��n4�P,���K���+�*�<+�NoFx��L�G��3K���F�T-f3*��-7zuM�C�M��4u"��F�}�xo��� �S��2�Z87�,��{$A�|.��d�X5��]��e�.��#7�/�����Z�q�#�b	z���$�tH��p�{�u��pp#'2K��%�8�o�<��*�k1��>ZO��v*��a�:�j[J��5�P��] V+xD�tun�J0�Ȇ|
dt]�%���-�ϱc�i�i0z�6�$ �U̺6@J��F�:H��Ǟ!h^�}����Q�"��L@{��lqm[�y᯹���s׭|���[y��y�y��_������z�����^�ȳ!�?�9�S������짮�VmN&'��w��h�S���[�t��K�+}�ǹG��U 8�O���m�W��n�U9r��Ǳ����'���e�޸��Q]ψ��`��a��*��p��ZnhRb�Y��~.�@6��X	�v�e|xK6��Ř�����
!�p�(U��
�$~�G�J��O� #�:� 
�J�6�;-�U{(�<|�\��)c�%M�s�(k[f���Ր-�f��Q��,k���3�K�p�L5h������ODhneCF�����Ri����ޫsQr�D�A� ���(�v���	Hсd��Ji���70�ݞ㑈M�V7cu�P	�Z[����k��i�\����C	���,VU:�ߓQ���jJi���Ć�Ԩb�����;�W���X~��?���d��ĨT/-�؞1�_��)��cB�"5�D����)����ҴhltLV7�^m1�whvL$�X�q5S������K�<?���½č�(0o�L��x`�#��Y����vJÉt��ǬO� ��J;�zM��3	�i�5]���B�
���\�I�?q0��7�5��J�NSȂ�|0��q ��!�̭�m$��[��R���O�B{f�S���0ֽ�Ӥ(#�Q�v����ߑ�<���m��Ѥ��-�WV�M�b�f������s�˙�dB��ݘGlu,������ bi���(4P�Cژ���ٴ���p7�^O�l�I�B��4�lH�� ';X)I���'q
-�HD��a5V�����/�W��~�d��	Y�/Ka�%��էej��,/��܍�y�;т@��_���R�.�����#���<&��m�q۬�-���~7�PȽ��9N����~Y�X�յ�ꪫ��|(W���޻� �����Bf����JX9b�ƻ�i����ֆy?4�{���˨@Lɋ'���+���Mw�������^�@�+T���$���X��j�a�N{}�0���V	[��p������\9��O,����_���+H��O�:�Fh\�V'd�L��샇��SϽ.�ʠ5M�y)�r���k�=�htcc���A}h�ãU&��d��������F��Q�.Q0 ��?�׎l���:��1s`mҗ� �4�N��H,ml6��d�'�/pƍu5��ձ�y� ;l
 �HZ%W�}hAJL/X�V�W5[ј���puL��Ɵ��6�W�f/ʱ�o���_�C����͐/j{R,��[ �d@��T�]��)r}B婥����FR$��ۤ��x�J�D�R��u�-�s,t��&�2y+g4[m:�|6G���U����� g�9��0 �v����ȩ��Lq��m�0��	����ӀG��1r�g�����Y�v�a>`ď�Ub���";^N�ވƼ$其D��$��8Z�cs.,��ɍP;<�q��q��ps"��g�$pS�B7���U���SB�����g���?��v��3i88pd���#^�g�U��ZF�=�n2}J�Z�n�F]�P�4X�sF9�j�>k�S*�3�{�<1Շ�,q�Q���\(cn6�sƭMl-V�8��_�?�㿗����?�ڏ�G?�I���~I�����X���>����3��vЌ�%�O�vu�ׁ~X6(H&��ޔ�sg�����;��_n6k����@9�nNʅ���N*��xT�juKJ�!q�kY]X��x@�7Z�uNc� 0���8��o0"[�C+��7�ɭw�&Ս-��ƃ4ܿ����蜯<vJn�rD�砜xyV�yB�_���rW2$Q&/�nM�aE�F��@q�_A=<���5:B����P�a�59����5mا�y}
�<x�����Jqaj�Z��V����e���kezf���B~�����<��]sX�����!K������c��k����uyM��Ê�jd�MP>4I����g�
����#v��e&wy�G�c���XY �AӖz28��k�x�n:4!6۬s���6�M�N��1=w�₱���u�O/�/ʓO>'�]���0'��-]Ù�i�YF�����v��冽�L!�g�$[��~�yS1� E`����kM)V��s�&���^�*��t�w7�X��,�+���p"`n�����tz=7�cv���+p��0v��S����=2a���J���Ǝ!D�Y�/&�OȈ���QYQ��QL����OҦ�8('E<�5@�����i���T�~�i9b*a���0%W�Q� �oMO�qN,I�F�g�KlDb}<G�ixy{�����-2�?�12==7Xp^��D\�#���dq��1��	-�B��J=����X����"��S�E�IZ�M�2���:�����([S�]Ϻ�=_�Šl��)���R���F��@��܌��]=�M�#> ��k^��C��/��/|~Q�sNJ#�,.�4�-�g"\]����q�`�~�Ur�܆�rX�ͪ�|�Mp�#$b/��\Σ�Ee �2$zy�����i�pǝGei���yI�/Ϲ���eJN�h8{o�Ay*7_�\}Ť�y���|��#�ʸ~�w����������Ծay����S?�=�_�����eT�Bሔ;M������/X�Lb؋-dn�����1�c��7<5`�¯?�(Wۖ7�s�|�k/ȗ��������޻��M���-�=,����/�poln�ˤ��q`��~��V�R�W����[ZC�eB^|���lPaj�u&�����t�'AsS��'�� v�Z�)��B�]�̒��AbY�e�ܸ�xU�gLӦ���k6�(JYOT)גŕ.Ǩn�	�D3��s��326��<�?��+R�u}��kee�2��WVCX���@u/��H3!���^U�X���n��p�Ȟ�F~��!�1�$�.� ���ςa�f`Ki��g��?�3f#��Df���^7��ݱ��X��Ŭ)�W[?�р�Ei3px픃9�f�"m�"�-"���0ؖ8c싞�RE�_�:}G;�2K���X�~#g���;�qq�;�5�c��;���C�6��oMH���dd$#���l��es
F86����E�>-&�Ewb����o�t!�K��]����x�/#�w�n��xv�RN���Q�|�p�@� s(��ּR.��P����;����(ϧ�N�eo��ϝ�l$)}+��Z��CF$)A��p����哿�'�������ZW��5Կ�}7��vU&�UF���Pr��7��~�Ey��R��z)Xӗ���ⶼ�יA� �T�Z{�b.��c�-���3)$�����AS6J��7}R^}}V^?�v 7����b?3J�N�l��;F8�Y��B���ڿ�'.�Ȱ޳~�}wTdj�y;X����׌���#��}w�h�"���㲿;�uT
�#�XM�%�S;�+��������}�&���[ؒǞ|�������WOΪ����k����>iIJ�AHB�8���@ň����۳OS쒬�7���^W���TS���)�`�BD�3��8�we�>726b���;�Vbd�Ɵ�N*�f�0Q��W���
qmo�Cڮ��/I4e�p�n�f�Z�Zm��MuDC�R��k��V�kEV��W���e3�(�#��s��b�0>X4e*�9���R�NrB�)�T6EѸ&!׋j%q�9t�o���2*�^F��(ѩ�%��hRG>f�.��z3�j�v�xELe�|#I���9x#i#���������&D�;��� ^��r��)�5� Jh�'���Y�x�hK���
|���ZL�I��ɖ��{��G�Z���H����/=F��`FH���NT]O:��G>��zM�e�@q����G�ʡ?"��0�b�ɢf�L2�Qt=�frA�ҋl�1DDm̮�_p��a����u���U��yn��
�-�_p�+�`_44��=;�U���h����U3Я��*7��<������馼��_��������G���ȭ7^!j�;���\\��զf�z�a��g&���{nȯ�ʧ�{��{?�~�\�uj<Ɯl�VtͲ=��c���P|�^Q���M4��\=&O��*��`*ΩQoǕ�b�Sc��tI�<< o~�ay׷L1c��#��vt�{��Rd�_�;B�:8����rӈ^۽��?��b
@3|�z.���&��xH�K�ڎ��^ϸ�{j��`��q�0�[��?�YS_]ۖ7>p�Ԛ]�V7�t�<�ܳr��R�о�+����jC&��=��Hnb�!}�]u9�����;0Y~��",,�4uS�tc�,i�����P����!}$K����i��6p�9�J K�%&�k�we��-��F8"xUnࡁ}r��9~dAh�<����T.\���G�ʓO�Jp��9wq���-�0�h�]��E����v��b�5D��r�P��f}+��W�m�F\4�u�o��Gyb�&a\�n���&4 �-��8�oP����*'��5�Lri�ͨ5J�!�k3�k��pu^��eR([a�V�C�c9�ufϢ�t��?�8�@RaAN̊!8ҋM�kޜu�4�5����[[4�Q�Y�����(9�-�g5bc��qo��Bt��8��JR\/�Ϯ����w��;�&.���3�t���Dx�ˢ�6���l�[&�����0ŕd�CB�g)t�#��L�x��)��s\�5��.{cf��r��"���M�����؂t�A~&��B,?���.=r�K?�)��O�Of�o�/��G����p�C����K��U}OY�ͬ�N�˱k�z�Ge���h��7@�yfʝ�uM�N�l2r�їʀ/S��䙧�����uu�%J8_p����K�ܔ�Ʋ��_�^�u�ڎHdt��-��S�&���8K�E1�]S�P�������\��?,�����㋲��-K�CCO61N��YgW��c���do*�`/^G�W��gΰL�h�*G������\y��n�H&����w��ȗ��"��� �F{nvU6Y9|`T{��=4&�������$u"ä�'D���ab@j��(ȸ ����;�jFO��.�-R����(�I�cj���,�pHw�W�Re��Kkl`Şe
ҕҨ~C7ʺ:���F��,(\5����o3��7 �զ�2��s�Y�n �{ހD����Rº����X�hI7B�k�[Fm�΂35�`�VK_�R��Ty;e����=�)��ݓz(��R���	JHZa�Y�NI���W�ǋ��])xZg7д��6��r�0=g-��g��E�6�ʅg�QcZ�G�,I.o�^�.��[&0un�l���}�>��ס��d%�kIi�'���vѳ�a��Cb�괺@8']=Ⱥ5�L�:�u�D� �P��?��m:R�fo՚tn`D�i�r����9��{4��gE�>ىg.�w���l�* ���Ѹ��)����3W�g&	^P�nn�j`S���U���R,edt�����|����c{����X��|ǻ�/�|���3�$	�|���0x8�&U1�5�똛��נ�	~�
��aV?�;�G4P'G>p�_��	y�1��O���B�8	%�H���WE��KqN4@ܚ?)�z����dtė�S��?�T�IG�N\u�ҰM?6u�J9ˠܐ��j��$�ݷ���ٔ���T*�|�R�U��}l��|�� ��c�)�(dZ�&�C�J�ϫ�d`�lo��f�-O�0�ƫ�zUV�_��J��>�:�m7�N,�~�\ifP�ddN�ܲ~�ڒ�ͬK���������!I��h���-`dS�� Fש�p���C�Uc$����iD:�>ϠC���F(6��9��tLd\��w�q,=q�>�%*��ɇ5
DQ����Ҧn��O��|H���p����F����!I�C���Z�'���06
& ��H+�c���+�]tSh���;����l��Ď�\%�&�R3fe�|<�B��N\m�g����.����ˣ�O	���Y�V�i{l�4�2�S��1q��U3����n=��ӯuӢ�7_v�9��Ѯ���j[�$�8P�4���}�����}1  ZX��m�9����Guo4b`�����z��&�ٵ��6f��ad�)���k|��y�s^?���� ��E.7���XN����H�"{�{�y���H��m�r{�ow�=w�ۻ4"(�LU�J-Y���^.�[�ӯ��m��ÇG�������}���ɫ���&������enaE�꜈<����4(�mU�G�n���C�W�]df248���2�V�nN;?�F㙲�'�9>������П��f����B��΢:kF�n�g�������< ���H@:-��w�ݥ�e�^��o��N2|F�6�!�����L��1?�ן��_��/ۅq��C%G���c�[���"PD�()�� �:�$��b]w`h�
��Mt�-/���jM^{}�6�n�/?�(y�z���n����mK�ѓ�z�#�5e�Fqۈ@�T�
7&v@���JVg��w���?4���Mx��&7�����<1u�_z�b��#�Ǆ�a�҄!���P��׈������4��V���E>�� ��)�:2u��bE�"�a@z�-�����p*"�~$�ڭ�$`ڻD_`'�l�Q�;�a{ݲ����ݣ�,N}�5�`�[�4f+��ia������Y"����I�*B�4��pה�ww�!���:�e����:��,�G��T�������#��@O� ~	nF|f�ҁ����|�$��wZ:�������b��e�O!^�)�H�Y��;�05|����s�ĕ��Mg+~���q<)^)�&���R�t)�n-ԶLLܭS@��,���� ���)����s��]���Ib,�%��@�[�˲����>G6�&�,r�{�	�����3fǕŋ��H��~��o��oU��_������g>,�Om�����Co|�����oy�?3����4K��p��\�]w��c�����<��5�o��Q/j��L�l4���ё	Y�mKc�+{�rr�Y�5�32��<"�8+[�tL�;��5;3RW��h���w����� ���kI��F�uϯ��k�� L1��������^��������)ёxc��[.�>J�8����^��O� XB�����[)��`z���$E���hLm�Z��-Q���p���ꍂb���$�z'O/s($��E�T�� Bܨ���i�� �:_cmo�a�#;lT{�Q�bzo���0CY ����$���2�U*�V�N��3>N�e��NK?=6 QF��=���2�ͱ��H�q��p�h|@��7�f�`{�F�CC������/���C�^�J5B��ǌ�,a�bD�`����������j�0"���"t@�ҊB���܈�#�>J$���X�@!]�\��w��)R�1Y�(�d
��wG����N�=-�f��݈��^ ���ގq ��­O�rl�A��̓�D�R�@8�B��Lq��r��AI.+	�3lX��3�N���P2nJ��t� A���~Ĳ��"f>�^l�M�������~����i�r4Z6�ș�Ӡ`x��,�T���������>N��?F�V���(��D�5$��n�8�K�OJ�i�����~�`��k+���"{���s/�$?�#�-_������iy�ѓ�-�Z~���| SE~�?��ϯ�����s�hԺ�Ī	���-���m��uW>�WOK��#��$������ێɡØ<LdttB`������G�̫kzfs�����2X
e~K�Ґ���w�(5"�7��kn
lie]��F١8��)��������x��RBЈA��*���E��ʸ<��K2R���Z���j�P���E�?�Y�&Cd{u$@ߌb�zj�@fU�M��n���zPs� "�����a~H3��`
�l�d�j��M#6�W#_҇\�o�<�Ѻ��i$U�mJ[Ij�%p�V��u^1��#���1���.���6L�:jzmy".��g�s��8�f���1�O#>�1�)�G֋+Ly�NSwP�g[��1�WJ�G������}������M�-��eF���f<4���H	��\1g�4���RX*K��@��G�U��`/��~���i:�lt�C\�.���{#c{���:��W����u�F�>.����!�]K�ؼ�ƒN�A���F\/��΀Ɖ���~��
C��@ܿg?U�N��f����v��IL)���|t�&t�8{$�����hk���?��<��VWL���(�̡;�"�5!�B��l�y�l�ᨯ���Glm�>���`��=����v�zw;L#���]P����c�����Nى�h���������� ��.zL������Q9~��o���|�o��'�mo��O���]��:�ɽ9�?V����'�g�?�q͸�7�;��1��͖X#� �Ы]^����/�H.���u����k�;"�]w@�~�9)�ȩ��������[��r��=��K��ՅځL��<5�a���n�g~�����\{�7��?�aӚ[�u��Qt{�Er9?�S��� �K[2�oL����C���A�W�Ҡ�F�y���"h�V�ܳfY��]T;j��������Rv�c��r]���h��!a�Gi�aԄ@* b�±6�0���ĺ���+�G9
`_TԀ�-�l��i�pʾ>�9�!�9F�$�� �8�^d��IzJI0G8p� �cJ.4'�&d����ي�����[����!�tC�W�,[�ɑ]��N����V̈��o$��!�&̙��q����}N�ׯ�u�oZ�d5��7F�x�h>'���3��m���';���
<'"����hL�Q��u�|�NOr����&��~T��g$tS�;T�I�d#�jHs�4���Z 1$I�0'&���j}��額�^3Ҥ�{���C��k�9��h����A\�K�+l�Y���Ҁ�#���PO��5�����MJ8r�`�Ku!�� &�9���~m=}��~ڝm}���uN�[�h���G<�)���`���рXoh�N|k}���w��^<w��wϝrxr�e���~�w�7�,����$?���Z3���u�3�\C����䠗ڭQ����ť�|�Ϟ��_�J����������xJ�RGf.l�V���eb�(O=�@�=ܡ���ݏ��z�S*�0ސ��/���SV8C<7��Y��O�ʿf��IF���x4��$6���mݧ��>�mo׆��G���'d�Y�28�a�m���	KÄ����'��7���%�,��{��[�Q���g䊅A���PC�U��Y@�<��`^|��e�d;��Qb�R��� dˑ�N�����`/M������6�<���� �d<ِߟ��a�0uG��>��/I����\�mh��R���b�qtD6���賋@� LZ�R�d��"���}bBA ��=��ܪ��K�9��T�'�}F��1�K	IZ|�'��(t�Ŗ����@�����9=�0���!���.�{�4y&H�{��!�J~[�%�0���`��}ϡ6����N�ʴAPZº���E&�.��Z��3zX�4|m��ՌZ�9�t�|wM0�qh�����>��&�`ٟ=��d����dc}P�;a�P:̄�����sӲg�(Q%x4/�5#�b�E��1'P���E5Be"[�zn4k�6�rdK�^�?G_�]��﷿g$m��5vF��O.7�;�Gѩ83��<7:+��zqQ�����W5��ҩ����>�>�_���܉�˩S�w<̟���}]�`oHn�ji��
��"��C�h>'����٠V{I��V�L����}^�-əs	{e]3u��,�4$S�����ِ�\��n�!�k�m��׭�dz�.W/�-�:�Ŏ�/.�ĞqY^Z�0�g�384F0�����l������ߜ����pi���^�����}~�}W��s�r�ަ�p)�v�gsl~Lta��O?쑔M9��������P�Z%� E�lL�_/,b]B�]�3������8���!��1�&6����j4W�w��CǱ}C���l�t�w����Z9��N
�"+k��n��&�y�r��	T��-څ����0��s" ��ێ	)�mp<{]F��l�k�'�~�0���H&���e8$���Ǡ�_�l�;2
U��MNR�1�2��(8>�e��8rS�!K[F�� ��*����Y�FݳF��U�C��K3/wQ~�8�^���L�ѩD��S��$�mͮ2
kԱ���1�V7N#�Ty%۶ �^)MiXc�Y����,��Ti�\q{/`���'�s]l�� �����P7��麢1����{� 5ņ�Tt*zȇ��S�5�:�t���s���xqF�~��Ǟ��x�фo�6Ed�䕖zA�z��E��������� ~�wy�pY���)�g_kk[29�_榫��?�?�o>�A��W�w�[�u���*��^Ǌr��7�h��(�������Q딄-��u!��$t;5'���L�4P��{]c�h�>X�}8�?ۖs�y��d=���A��$�G��!�ą�L�ѲW]��������;�CKV��Q��ꝁ'S�IY3��ՃN������{&d}u]F v�i���Y�W{�7���A���|�9��M99R$L�`�ah%K� ���PV����4�Hʵ��Y�X�,����C�V#�����Z�M)��A֦�O�z�lմ��������bu�F���""�&`�V�Fjq�d��di��_��cj\�gX�t.!|+��Ʀ��rm��M���������%���jM�&@M��\�g��%.�
Դ�H=���x�zs'�]�jZ�!����[V��z&��\�1vM��w*\xr�8f�ɗS�z_~�z�mK~y�3��h;���u�2�����z�(آ&αz��Gl���i�xW�_���;î�"vMc��%�3�ρWwW�k8v�J%�k��52	����I�&(��?�a�"�ó¢2+����Ȓv�FREA*������'���ɹ�穩���EMF�1C06�����y�%�\����S�u�ގcyLeĐ��k�>? ���(xw��/����3���b��9�������J�)j�[�j�~��ӯZ�`0ז��(�����������ğ�K/�*��և�<('^�(7�zH~�?���b}V���y�9���5�f�2��Au(WfY�� rЁ��N飲k�#���H2�oM����ɨI��]�*d�=����tk{Q����-�B-;N�}�,�ogff��4B�3@���b�	&��p��Cj3ԁ��f�/��I��c���1=:*��������;!TÛ!��q
�Ef����B�25uP�Ą��b�?pRv����
F����C�n��R1���I�%��Nz( ���f�,j�|��t�Ǧ*�'][ݔ��,�i�.��$�|~����R�5��X$����W���櫫�N_��^��O�,��s��G\шhx����Ե7�m�n�46.�9�[�R�HUrD@��� �E����>�����[M�m~iC�F��6Zl��w������@-[+�栁=b����)�21�gwLı�Ji�[e/D�XkdD��CYB�>w��K�F�-'�:k�����v�����C����6�ym��w���4%�m�3��1��f�8��9Qd�:�zD"e+�|b'�OG�-N��DP=�����:8 TSl"�3�(ԡ#��K����3WHb�a��=���K�^�)h�j���B���fU#���e��<0)�?_o��Y�	�o������<$�f�I�� �0��
���>]�bkY"8�]��eYU]j�ck;PZP�@�Q�"`dIHH��n�;�{��S�ַ��O�>xs�=������ַֻ������+��'�<,g|H�_s��~�i5�;Cw�*���LyBu2'}P?s[�k��-[[��UＴ
k)�J�������gc��"_����8���S�obp�����$)%C�����|�#Rs1�0��_�i��uފ�&�XN�M {�a�P�Y��hsm��m>	Z��C��9���5]��=��P)���?А�|�K��o������`�@L�J����5��nkL��X����K$�Nlo1��Z�v�>�^�#ǎZ����|U|�%��i���^���/H�X�UG��u�2����\'ݥ�i�BOݖ�G[��*UTFre>8��,1�U8X���|��`S�J���1�mAQ(1���ލM�^cX��vqc��j�=�"'���J��8�(E��P���1���O�<�7���4���׿�߿��-�� ��x���S���h7������ׄ,�̙����+��@�u�:�	~�H�ꘃ)�VD3do�6|�^�Y����ɡ�|�2�_���¨c�m�jB��\���"DVZD�T�����}HqI�}z��{	�� �Mm��p��s/|p��A6�b|����Oՙt��M�,ˌ�Qo�y���=Dޘr��d��[��?\rm�Q�@��X�VqH6؈.�<&��Ģ8��F�΀Ar��W���A��:��~S<���G��m����!4��r��1V|"u��+|2�y���d���v�̆��تa���a�����|S�z�b�ZG(*����ʎ	�0/U�1s��-���#�,��M��H;g�^\� ��3�g���w�������Eo�WCSpr���o�İwU� ���L���ۻ=o�����Vei̱�f��W��dW�f��ƌIӽ��Vd�l4�o�鐼���5�ѡD� ض��\:rn��
J�yx��d�R�Ά��_����`�?����Ăs�%]����<������Wd�e�mIp�-��-|�^���5ǎ�������1f��f8�I�Km$��*��*+��o��<r�1�w�Q�>~P�gч�$Ji����N:�.��'�<'�����N�6��>8;&^��Q/�����7}�МѦ�a���D���*괳��Lh�g�W_8$���|F��PΛ�n@�{����*�wa{S:~#A1S�,�]d��&�gG&%�r��S>�3`oo����&��u�[f&&b��лu9W�ב$�9��6�b������LF�����c��7/���`
�����)�;�|��LJ���E
*B�xƞ�ʱZ��^�f���j%���b>s׏��A��F��H@�2�׺ ���; ���P��
�2&���^dՉ��B5_xXơ�SF��qݣ��fh��z"l��>�oQߧь}²!������%�i*Ϲ�����L:6���J��� �o}�r�`mw2�(���W˰:�y0��L*U[�eX�j�"Ѻ0f��u�<�ȣ~����W>[~���\~��#?��.���{s�ʅH���?�-A�{ū~���+�1�V�C�3�];�р0��T'��3+��[��V�0��O�"��	l��-��`�Ɉ`<�a�������&i�����qve)2�?����@n$m���C��W~�P>��� auII�O"�nteiq�I����R+���`�<{�0fͮ$3��>�.��ƚ�����d�qA�}꘾��Y� ��� i��2.��L	SV1�9���J� "+W�:�7EF�����Muа�gA
��(!WP��z�C�"� :�����2�%
�[��,�T1+2QJ>m~E*�Y�x���+}������4���Z�0:�pQV��x0X�8@��.u����;�&���r�ѧ��t����:�0L��PQ)����p`%��@B���O��r���Ҫ2V�)�\�~�YS ��_.0AgP�K�rߗ��,�[�L�8���ʺ�av�6|"����.��cB37��a:Q��[/DW.�U��N�i�0hh!Z2�i�������k�<1�LYVX;�mQT?�,���
��x	�4��"����}���\�1ި�ۍ��`�['w�sB�h�3��������餣2��jS�)z�c�R�@���nu�V�W�bސ*�Ϧ�g��m��!�\Ӎp� $���Z�Y�W���ѱZ�m��	��>uy�|���C���������G�{xP�?!�'�g��Ly�u����S��o~Xv�~��'`~� ����e���MH�mfK~�mH#�`_�j���|�2�U?�ݣ���v��2���=lŜF�1��d2��Lf�>��D�n.��]�����D��;OU�r���k=_=_ܵ�� ]|�_��X�Z�0�MAW5G^~\��9���ZS.;�,��I��d�?��[�\�͸ɒ��ظ;q�\ܔq�I����֖}�C*l��1=�C���yqK�C-�)�sİߗ����8���r�g�,����d�аld0�Y,�Cn^����d��hF۩<�ϬU��ʥ�8ȁFf��:籼X�����%����n��}�ak��g��9�&�}��#\�)+���ZM`�J�G�!7�j��8z�kAt�g��0��#�'r $cp	��P$C�\ �l�����Ɛ!��,,��=� D�IQ��w$bq��Ťa�Y'��&E4-�Y"���²℻�����j2��h��0D��=U���=N�̈�������H)+M][��ב�EEt�Ȫ5gf�I7K���P��i���b=Ѧ$�=(�T'���{�Jp�E��aL9���2SG�V�l��
⫘N1	�6��0�1��,k�����܀ q�ᚇÑ,,��0����6}N�`��W'#(b�-�Kz/�{R�!l,x�ީ>��$Yt�!<�SK�i��Z�ħ&�%��:�L���+F_���r������~�M�+��C��<%?�#��A�̙G�^�Jy��^!�yQ}�%c�o�I��P�kX~��)�-u�X6|�2�s�����O|.�=��3r�-'�-���p�	YX>(�K���m���k���m���Ij���M��_���e�b!�D2�𹻍�Lx����V� \' ���u�Ǆ�����$6��*7�������C�~� ʑxr���o����H����A����r����`�����Yd��@�{�l���c�������a����*�������gp @����~ED�fN0����VV�Wr�s��RPޣL��*�6��a�t�����%,*���t`� [a3����?Y����|���ɣ���}<������`z|�Ȗ�\��J"q*��3d��y������3Jl�qS������C��t��	�������X�Yu��5��_�:�>f���ƗS�'��Q��!I� %:���D�#��#e��*���L��ި�vOQ�-����<�:)mЧ,�@�3�X��bBp#rL�-lDv�?ie����t�Ѽ/����%'�r>��T(�m���8
Vh��Q�F�6��Мj�9ke�Q�����S���٬�V& i�Tl�
�`d�O|G^L�ό�
��
f�S� ���0�E�� ��*;��݁_o�;os�}��W�
��N���������U��UԦ��Es��i�IN�,���|�����_�W������:����?��]�o����W���{Qȯ߷-םZ�w�ܛ������7K����.C}e�BhJ6���߷�;�=>,��[���_~Dn{�q�d0l�O������Srn}���^�%>�#	G���}Bn�ή�oNe{��\}�ъީeJ�x�?�a.B�c
�eL���h4}���I������{2�0w�?����假��KN�8���ē򤆙���:�A^v�*�l��g�͵5z��H��͘����D6�t�v�E�AN�R�$;>p�z��#3��ޘ%� �����~�g�=����B�B�K�`�����>��UfQ�����P�� AKʌ���h�Y���=x� 3*(�9`H�&�p�w���&��)�naIEfGb:F«��e�Xh�u��_`h�~D�=� ��XO�fG�w>PP"}v5����h9�����Ih��,:�{J������;,��;���E4H�JME�'�K��0�dQ�.pF�3�@3H�M$՚��V�L4��8�U�,���i�Kr�vı6�����@bq�c�T�~��1J��ډ1A���lc���|g3���Ӂ<[@R���}����mLS@���j��;��C�<�W��ը�7M\o
�W�*�{���
����k�?A_����ɐ�!�Se�N��� �A���z��_���;W�]�9�
+�מ_�-���S�����!H�'�*m��{aڭ�Ǟ��Ə�����0�bݬ��u�-"/��V��G�J폴��VB����&[0�����Y,*���ʚ��/�o{vK��ңr��7ʗ�~T���tҗ��������+���i��6F�IA!�WZВk�jx6��~�>#7�t5N�	�cT�Yc��oQ�� <`�X�f*��MSc����l��-fE�=q@��В/=�+�xY򑿞�G�N3��vw�-�ߣ�G��՛o�>|B
���f��?ra�LK��(���`�nJp�F�����Ȏ1)����m����}����U�6g�@|���G�q�0��Dm����D�d���Nj֒�mw�@@�fPJ����0��~���f�&8�3�L��U#�3�fx�o[Il
��'�ڐ*��[j3Y���L�Q}p�@��8ٖ%<�����4���6|&X��NE��]�,	~���`�b�AhD	/*�5Ѻ��^����7 ��	N*B�0Qˈ+��ζ�4Hx��J�MC�S�z��fw
�8:��3%�rlӬ��;�'r�yT8
�U�J�U�އ�������<m���Պ!R�G���c����9��;�U��7�J�҄�r��7f�G��+�,*���5�y6�3L~Z�V���Ly�K��@��yX&�"�@K(̕�=
���2
��ظ7e5]>q5��k��K�eT�S{�~�ɼ(��-iF\��������������Y����Y��y��N^�]��w��/��~��ww~N��}���?~OVW[���U~��Z:td����F�x�.[ۏ��S��:�,��[o���=E)�ݟ�W���������o������&�}��o��n9rpQ?�,�J�M*W�����p�/�d�ڒ�93�׽�
;sض���M"fNR�Rݡ���Hڦ�����,��$o�dS�3w> Ͻ��[�I��(��&�`�9M��Z�+�=��R�ey� �v�����3������[3�Κ}x�3ʦF� ��u�FS�>pcQDk^v	϶��0(/�&�+��@��L�����x�E�ri����+�f4���9��J��Yw=� 6���YZlUY8���>>����o���� "XL�{��3�0��C��n�S�.�S��h�
��&����{l������+I����f� ~oʬ#���O�V�:�nvɃ:b3K�V�0]G�(�T �A����8�IZ��5s�Ձ�m���P��-/O�T~�L.���R[&'�kA�4��Kg�P$�N���vi*PT�L����Y��Y[�Ȳ�lQ�a#*�P�)P���Q%�@粢���B?EZ��Y|=���*ѯpj�h˹ �V��Z=�ϸ���91�ogEq��F�mMۢp�Y8�RVO�R��y�E�����p��_M\�t3Vq9���1����ž:��y�3��~�g��_�7�����ۮ������o����?%�3�w���H���W���N�8�ȅ'����^!�1���5]������aYZړ7��M���9�@��<�[��s�?��y�!����s��׿�6~�o�M^����W���e�e{	SC�]�:��m�xW,ʬ8(��En��'����������	��"���}>�64k�<�h.q���h`"6@U0	3��J���/�V>���}wmI�=!�����$�g�(x���i�՗�~� �EZ��`:P�+L����FT�H��l� -2�*>�&���	>9f�� Ѽ(uP�����aYJ�1~2�0iN��Uo:܃�e�����&y����:�P!�UԲ�@M�c�YpK�d��M9ظŀO�'�m��ҩ�zê
J`�����ZfsM	8���µkE;5i�=ӑc4<�¦�5���ݝ*�Y�1�dF	��\<d
�����E�!f���#�pP�ZB@��^c܆A,jH[�	A5b�)`Eh���~�*D��w̵��ލ���<�Z�(�
3�Y��~\�\4l6D��i������)97��F�hT:q1[ԟ	h�N���5؀(�<��?r�]��6GH�|�3��:���1�Bk�;�̀J����fO��a.��E�����N���XdN�*��Od4��	KS}�� MWV�!���Q$�;ӡ���ԟ�ţfb�sT���(	C�iaoeQҝu~����Oy�����^�����]���N?x^vw��_�˭ϻ[O6������_}�	_Q4��`,}JvN����i����'*x��O�����`p�,���u��Y�u9q�zvg6�����~�����e��>�l.�����d\ͨ
P�./^�?�-y�{>/?��
�8�0J��1�ܤ����Yl�:KH3��2.lQ���ȝ����s�<���G�����q�=�����;,d�����}!�X%E���S����_e�.��Ƀv@)�C�h$�7q�%�,��ˬd�'�6���O(6x2Z"���C�IaSK����tb�fb���Ҋ+��t]&��m�H.	�TT<�R"�B��8����ƋuЃ���C�<tp�LGc�2@����K���Fh�h�3��.A� �o���+%?ۑ�y:	��	f��6�N0��!G9Ld���Y�k�*��Qc`fں�������h6@Ƅ��t\�R�MM�{4�UA"��h��5'(
��{�;Ί*D#����k��-1��"���J7Lmm�����Y���-�]�F����xaZ��~��ޖ�qF6�W872�d&.˗`T���	M��A��*:� D��n��ʍ.��%O�������
`�Oc���@e�/�DH�z�ޙAΕ;��Q$��Q}��Yl-�ޔ	�K�7��Ō>͑�CG����uox�@���NV�o>������}�c�s��k2���ٷ^ŀ��=Bq�\��J�C?��)����}�c�����g>wn���?q�� xu�0o�(����������������#>h�5H ��@�dS�L�-�d?��lI���Y��pc���X)M�5m�C��� ��(h��S9}z(�\��3g�>�İ��v>�AW�}JL[�XP�#���L���7��u����?��3-S�sՔ��\/PԐM�8�[�#glF6󑲙̔��l"����56=�%�HЩO:�.J�f������S.��G@��3�H�l)a���r����VB�>��*�WT�����p���=9�^�d}O�ծ�"p�oߚ:��F���@￯��sNl9��Kd5�힤��̢p���A��8�}#�m��Hl�-,�d��o���6Z6�����+�,�X��2�KkN�,�ltg�߲�<�%3H��S��!�r��S��a��L4)`��f�Y���1C�/���r��54�ݦb��i	#�ya���U�B!���L�ek}�ШsF����*�Ka�\3Tn��q��`�
�Ü�BK�6�:���Ƽ���WY�����l��Im��[יf:��aB!=��Ќl�9�O0�CE�3�C�`���9dÈX��fQi��*4�� ���ϴ�[��~E~�߾Vn�բ��fp����ɫ������^��&d��+�>S������-A���t���W����qO��m����YY�����.p_X\��a����j��xR9%�~��>���e:��AfYF>K���݉5�`�c�a���?�<�)����}G��0���s��+-@����V����=��Ş<�͡��oD�[��;��E�*����X��o��DI�(%
AS���q���>�_�S{E��?讏�1���*V�|ik僪�*�7�H���n)]D4����(\k ����z�Ê8߬�Θ�A�\L�1j\3�g_i�>�Bޠ���ř�8$��Z�]�,D���$�A/z�"����h�r����ل��0R?H�4����=�=f���	��A;˝�ȶnm��y=�L�[��SO7�����rR�&���B1��/�x��0gl�V:hlix�����c楕��T�0s��x74$q�5}�26(5L���qBa�ݕc���3<W����kt��q6�t�(��¡D�5s\ݠ.-H(>c��Nʚ���v��*?S6LDH�A�$1w��)ި��VI��Y^�a°z����k��S7�,fo��d�cm�j�A)����z��y���jrBb��I��`���p�79�^g�RJ4�z����ŧ����Y̽���c�����+���'�w����_�A�����Wi!ؤ(	�n���X6��'_�����w�'�04��,�?|Zͯ�T�<�?���?%����h��)��<'7�|H�6�r�uy䛚Ί'e��J�k�|!u2�|~�m,��rD^��7�_|�+��^)!|� ai�m7�>�?�p(u�\&���^��;��C�ɳS����]�=B�6fLL�Ps�J<&��Us�+K~!c&(�K;}3��Q��N��S��`�.`�x�'!4u1�װ�~&����2�hң�VS��	���G�����6Eq��yA�0bcO5�U��FH��R�ye�XZ�3�˫��_U�!�ѧ0�]�[@]�!�^�F�?D��� �_��*Mjn4h"v[m�R��:�d�p�L��!r�`<>?��A�����\`�0��|��x0�`,�H��[��oq��� ��$<��?�Ӓ�~S�jv4�u��0�p��bd���m-s<�xv�{��Ɨz�^S3w#��*�'��T2s��z��ck��G��=<S�F�� t0o�F7"����ԙ�q�Ss�皈U�<{����q�h��^D��p�"S��(05��h���,���	Epf����j<�0��UJ���a�5NT ���tz���h����;�qr��R)�Ҵ�C��>�K++9+�ņ�
��whw����@��xxA�����e=>����m7d2HĊ&y��L�w�_�8ҕ�����_����Y�L�3Y���3d�Me(o�_P�#�4�[�dք�ڠ���s��H#�$��Xҧ����LV&r��o�O�W���� ��%�lu*U�g	�7���і�H��C��d�=�����'�󓯔'���/>,_��!Y۷_n�������������G��/�}_�n1�1D��L0g/	�!�q��z�D�?�\��㞮��%����[2N{ }�9��$�'r�7g��,�ЗNb47�_ǆGO�iI�,TWat<,�!yއ;���"3Ɗ�э���hE�m�M�t��ZLaE�dd�x�ܳ���x�� �&��0t�N$X�'��ih��YZ�ƃ�\Љ��4��)Lr��,.z��S��;{R�8��fx�;Sq=��Y!�`_&�NK�Qz��d��o�̍{�v����Ax&�G�(��v�����13>�E�NoF�v*t����pI"(L;�Q�:�E��xJyb��Y /�n���F\ib�>cOH�tS�D&qZ5Q�a��QTn1�N[Θf�E�Z�p��tI]U�q�+fR�M�&!�x�?���+,6xK�bQAY�������F��
��2=�*��Ri����努_L�u݅d�6�Ps�Dº�,�K��L�1�	i���K�DnPu��EZ	Dv�5[Ġ1,�=�F����z��¹�;�~�;�+�������|��U/��|�K���_(����o��da��G�8-������?��򒗼\>����G ����c�3�-��~_�>%�VV�{��n���1Y���
a���(Q��?����'�U$�,Rn�g�x=�_��?�Te�w��Na@	��LV(���@�v�Y�ȭ�]&�g��nOc��H�L*_��{�ϻN���?�cO����A6l��v����G���6O�2q��������B�,��З�Ξ������[����,/.�z۝�?�>x%���7�l�z ~��})����Hڻ�CY^]�%Q���4>���L)lX�d��X��c}}Cέ����2���>x5!��^����*�9B\1�u�Q�+c �e`��]�r���%���w4��:Ed6US���Җ/��*�1���_�g2����M��yF�T�7Z�v�L���F��Qbf;��s��2�N�7�/@E����A���:)��pO��q/�M��)�ņ��q��/΁?��I������{����y6����f�ߒN�|�t���R�&�7�NapL�����[y�ͬ�/	��f�b�M���\D�u���ӕ:�/zk�x8@�Qk��*�Dk
��#EKI�p�������K��1!K^?�`�a���i�H3Röm�H�T���	^�.V�`}�IP�*L���1x��m�-~@t8����u?
Ӡ��B2��6��^�Â�'A���vQ���Yx�G�^7g7�|	�*�4����l,�Ï���J����3�;��^�����j���\;�$ǎ/3`�����"w��Sr`�{�%'���|�l/���-�ʗ?��O>����c6��5��(��Я��Ҁ����;&���3�u���/~Uc�|j(q�W�����S0�f%�������_�ƻ^���'��~�s9v,�G�M�h�J��������Ei��Ŀo�X[�>��w�v>1j��=֗���o����zu8'K]wL�������x]<��\v�l�r���U~=�Y6�ȉ	�gfV6���7�lާN����]Y��� .O"|�٫�N;� ���{��O�;G�<�pG{��p��?;� f�Lz�����:qf!�)]^�)���M�͌�%s��`6���Klz���O,�� �L��b�4h0�7���#�Wb�5�&�+�lw��c:��Ǚ,`��&;A�t��e;�I�<46;t!Z�e�`<`%��!r�3$���o�5�����S6Q#�~��<\�W�4��f�b��U|>|&�����N�SmT���~Xy�Z��-z�Y��z�Ny�j?�f޸�N�U0�P��	��R�mb���D�<�H嬨�F��l� ��� u-W�P6鐒�Z�$�֏�L�k3c`�(�1��cNh��~�8 ��&eڴ�/�Z����	��`��j�H�Cf���e��P}����� �X��| ��y�J�+�����MN>��O�JD'm�P
���n��1�����g�����ZO�E/}���8y�Q�ԩ�,t[r���f�o�U�v߽���~Z����d喸�Ǒ�MA��6���:)7�d��_���w���H�<i�m�uE���"0n:�]���|r�oy���ߩ�gbF*`/"��lBlL�ES#b=�)�x�����s�>a�ch��#�=w��|�#Q���QЙ1�1`'~���T��Ȏ8`�����1�*|��؈���y��#�T.\ܐ+.����x<��ǆ��t<�&��(�e�+O��a�K��;��Ȑ2AT�ސ�&���VU���Z]Z��L�x�)��ʓ2�N������ѧ��=L9"�P���Anq���j�-��<3� �L�4:`��R3��(UiM)�r	��6d�-�*uE���=Z�\�B7-��6�a��:�=�i#�*�,�/��taT꿾��>g�A����r�H"��xS���{4UK�^`� w�{M�p8W?4d}�񝋪�ȁ�K;�́�uP��[f��-�tI]�U�+OlX���ks���zG�a2Ն/���
�&6�+�_�l��ʡ�Y�dB0@�U;��o�!
^j%�2i�B_��`�P|�,�8Xf����Œ*xM���j��kLh)̚����R/sƕr��"�~Q����a�14!��nLd���h%Vȼf��N�jx4�ѳ�د���=2p ��Y���[����q8��+u8��������u���,����W�oV��L|Wӝ"Je�;�5_��Sw��/~�]�_���2m�x���Q`���2�\�;5@hv��.������y��O������H ��S����zy� �$������./H�g��p&�(���9���z(��	�4^t�� �7�H�E5A�uN.�k�W��$��Pth��f`�V�y�k_����)���F�P���kk�r��u	J=�٘��f�`ІPΡ�d� G/�ߔ�O]f�<�����<�fu���F�P�=,~�Q��v�>�
|�q��S��#qS����h|�ك]b@J�_e"4��r�!��\Q�=nh�I�i�#�$c���E����� ���FC�.��2�X文k:8��Y^'J�sq݀
YG�-#������&ɜ�S&@��Y���:#���B�Ѯ���Xȸ��C�`����l�d!Qa�ЏA�,D p�Ļ�0�R:c'��n�4��I��>�n�Qi�^�jڑM�`�U�kN8P#�ep=8K�s�:�oTY��tN���!�z�?�y����MT�}�
�8� H��Ǥ`⻊�`�f�#ꅭǘ��Am�p��YXv���s/M�ıj���\;��R�Џb��e���x�.<Oe*!�
=$dY>##
�`���\~Y��I����+��7�J>��_������{��:y��M��w�_~���+y����\s�Ay����l�T���>C-�HH(ˑ|���3h?���>�	_��@��do�׆K��vS�5�4���+z�����;�{���=������y3F��y^�����wj{'���-�|���	��xI��-�V|l�Up�3j�1�<`}b�Y�R�y�Q��E�8��$����,��]�?�o��ڢ����Հ �e��`yJobGvn:���5@F�m����/,��2�i�2����88� �Dy���	\�ȡ����rז�T��<񦣸��B}��Z�&l���g�4��eO�JC�͠�n(!�f�j��K�JR�����2�76��5��QU7p�$*3j��v���,hv�t�	|k��Ri3�l2"X�[g\�Sd ������b졠�|�Hl�꤯W�l
gң��62�}Ɉ�Z_dll>4^y�*���j��C�������\���3h�)IY�@�е0g�e�v���g��U�����dz�R�MX�0��}Ḥ��QC�:O���p��v��yO3�L+O�B������˼���D�t�=(/�V�'�Z&§� h����8y[V�r�qaا��;?�3w���e-ߋ��v�����*������<�m9�Z�w�����aA�x��˾E���˟+��'������;7����~y�͇�k_=�k�\~����&0�-V|��y�{>&?�o^����4��`�b�Lg���=�>֋O<��`��"�����[.�f�y:�4OB���+$�=P�_����3ur{����h㰿�(O�8����2M��W�U�l}���=�	'^Lޕ�"P���#G�C����>`��1��3����;Ų
�tn8������3eF@6���|�צ;����G�������hCa�mh�����9t�'QL����f���E� ���m�Q��X��f���l��(�s�'�VϪ�r�Ͻ�D�N�G�El�BUh5.J��gLA�8)-3w:�Y]?$l�I���Xs���VX�e��P�����=���[s�� '!N����@��X�S�A�^%��"�9Cg���Ln�Bn�Q�YS;�V/�pH�����f��aB�*�O8�l]��ޢ"�,G�5�`0�� ~�h3}^�i)f��.�l������3xy��*��5@&H��i�ϼ�N���i^U��f�4��:��,d�AcT٠f����,��҆s$���w���^y��+K���r��)���TrA5�;��l�a��_}�|�y�K��?����_�B��x�O��/��?��������;�Ǿ����W�R���k�̓>p7����$%}��>�9�݃r�O�]w����A�I�GU��M��0��A��b��n�K,��ux�#[��0D��7b26J� n�v8x�δ��<5�$�F#�༊�=��rL�4Q���%9���ظ��D:�:�!(�"4�a�1X��ޅ���f ��?���Vd{cW�h��l+w8=U8v��Ʌ,%��`Ma���hx�,3�P�c�f����p0O����"bAiT4!��c!�ǵ1s���K�L����,�E��
 �e�9�ͥ6p�"��VD*�
��$�uנ͑T�:p���2Xkq.d��u_��sA��B8��N�G|�}Ol�ebf!���sB<.�2(���]�K�w�y��uባz��x:b����)~�P ��S�!p������{!�t�/�E����s�+���m.�+Ğ����L�f�Zi��dY�5�R����G�=T��Vy���qB]���s�bb���@c�_t�1�G������Y˔C]�(��o��lmoq� {F`�U��DhuE��f�����LG�	��*x}2��ZA�6%&F��0hP��gQ�RX��l��Z}�^ߑ����������/�-���/��?�\~�ٸ0�o}�d0� ���G�:y�K/���-(n�8���_"��x��,kˇ>�)9pPc�������/��W����|V>����1m�P�������=`m=y�$V�Ow6E���Pd�u��ETZ�Uj#�U�XM��߉RB]2���1_w62�f'T%�ͭSX���Iq`��S&� ��[pcG�|c\ȡ�������V����:�����l:� n�OciX#��A���X��iYeI*u��B�n/���R����Ȫ&�*JU-���D�6��E��b��vq��ymF�
F�@@	
�7:��S)Q	%p�u�gX-7����S�.貆i���j��=]d4e�է�iZef��[��US_�J�~�0��Q�T
��i��I>�a�A���%�|.�i2xȚU#�Ł@��]�U�:��z窕���ƹ�������$�WYC$s�3ܿpuZ��FTue#/Mn4� ���C D�Qi�A�)�y�>�+����V�5h�`��N.|�8�6���\����| �/ӑ���]jk����1aa�¯4(k�9xH��H��b5���,-.V�:ޮ���{Vq�)�A+�W.�� ���Ը�T��^?�
��#V£�T�������?~T|�%л�����%�j���Z��W::�����:�4���+��|UM����>�G�-������S��o���گ}X^����3n>(ۛ������f!�����Geu�//(-��;K���^�q���7�(�l`�i�[�� �:2��EuǂA\�T�Ӓ��9��뻖��B�@8�ءO�q��M�v��x�:Jv�a'�$���U `�7H)��QG9N���q��������7iC�ܧ�v@��4SZ3/�p;4��mL2�2���!�� )E�P�r�[��:@�{v�?ˌ(�E��B�
�:�L�[O��2�K��B�4͍�,�e��R<-�gҘդ-��hh~�������������ߌ;'���1��4w��F�0���`�A��� ����=��C�%�E�EʂI����ZZc��O������wAm��!F�9�����UTY69����Y�6.;gS䒈`j�=#��;*2����D�`��Bʹ���Jﱫ �V#�*rSm���D��3	���@��ni�C(�z.��|�=��w�ve�e�`g�����,��;�O>��5wթ��=�V����Sy����"���kngw����RI�o��{�_�i@���}�����r�e�`Y��Y�3(���`.$���X>��O�ʾ���[��F�ģߏ���E�l<�q����_ܑ��o�	ݠxX�S�|�]}6)HȨ���ѷ�Wy�sO����<���~aK��������<&���/5���w�8��x�f�4V}��+�I��l$F��4T��JK��P3��a���{��cl��$��Y\��Ii[�=�B8l<cAyi������І���$�]ӊ^0�z��S@`��\R
��k��6�5e���=Iĝ�FgC�
�0�M�b-��uI�D�0,6t��o]h����D�1-�e��ޓ}��$�np�)T��Pa{��#e���m<`ѥa)�
@���t��KCCX��#�T}�fR��q��0qEe^K|���oݏ�ע��Z�΂�.�<#�b���L1Rh�,��
��]�@�/�6����1C��P�"��6d���TYSߔ�Q����~����|���� ��k�3�A@
������(a�7��RB���s���N=��ih�h�~}R�%�UX|���&��`W��򥑘Ԃ��W�
C7\�dw��RqH(�O�-�b|�=��{��ͼ��Bo�kR���������g�,g0�^��`��?d:����#��0����'dͦ���wu���>p/0@�J��x�Q�ԯ����0Ax>Za��n��|p�����^���XV�:����!/����$������J�ǆ���L�����$?��7�/���Io��u5).�g��vAz J�|��&�e���>"鬔{���|�w������ĉr�'�A^��g��s�r�����=�2�v���}uP�;l��g��M�SIgU�+��fHX3��	����!� ��G��g �K1�UI���!T��lG0`����f��!	4�,��2EÁ�w�>jv��F�Z͵nh��1p���yVR�Ta�
TPfӅ�d7���ёiЋ����H����B\���S?�WE��Xu�4c�6��ѝ���7f>(bHEG{�*�(,3Օ�7�q�f�t�ˢjb�S/e��ad��d Y�#XCŚj�����5��(����y%2������u�g�AS�ZE��r@4C�{��V�]��:�h��\k.��b��"c�D�%G�s�xj�ĳ�P���<���F��zLX$��da��Zm)M0����
y�����۰�D�_���X���h��pN*	�pHqX��L>L)0D76��*Jr������u�Cߔ��.?������@n{֭s,��sK���}^:-���'ϋo��%�nϟ9��٢Yv{��G����6i�`|-�,�~�A6�;�})������Z����J��\�NT�H9�q�����%tksӯ�����^/��+>���?/���|ǫ_���w}]~�������W��?���GO��qM��d��8UZ�T���t�L��Z�X0�(����j]y���f�D���O��v��7�I(��&���qX�-��jg0S,�)�����u��W�$g�B�̩s��Wj�����Ԋ��`��|�0u5�B�iw4��M&��$ӽ�33��yD-źR�b��B]HRh\<M��'��NM�i�Cc0��AZ,���TT����`l�m��<�9�n�Z�]�/�S"d�{�#���>8���fJ�_�f3�f��p�X��%�b���R��j���V+���&�Dɋ�����Ca ���22���x��m�>}Ъ�R����w���lZj�'O4�f�XS7��T8m�ʹ�O8-�-3�(��&�(xXlz��Fi������:�UÚ�vh1p�3
pŌ�F�A�N4�c��M��^b��ą�`P�ܴ�~e%uW����2ah��C��ѡ}t%����(��
)�L���Pu�	Bl,tȁZ�3�zq����us�@��M��}ޞ�U* ���:dr���O>!�|ի�3�f�1l�V�t	�p���9yέ��;���g��z���_��N?"��yJ�>y�ƃ���r�h���8��{�;�|g&��B�1蔀!���J��
������z���0���ڛ�����������dm�j��x�_���3���|�Nܕܴ��ݘ'T�-�4ZK>F���ٞ�'��|¾�|�Cw��}�M��X2���^@�����H�_��!�I�j�-��wL:�h��v�Hmsj�7�d���E@�s�����5@���FtOJ+�Q�5ʠ&tWIP.�t�i���~�2�E� � ��EyLd�m_�`�#Հ�Oƫ�i��)x�������`����b?&������t�/4�s30�F�fzg,��b1���qv��S�٠�l��D�����^�A,��Ӭ~��[	3�VK�|,�4�hsf��\ *L#��a��۪6�lC�)�^�F�˝B(Ҍ`���RLT�.��`L�قM����7�����KR��zC�sj[�)#�\.���S%��Ц���� ��4j�.GS�9�S�/%Q��g,����l6܅�=N �itDeY52]�%h�����X+� ���ߋ�e��v������Z�'�n�d�2�p
�Xu:�&��K�`��gS����=W�����cCZW^�[,�8�/��S��&��oM%$`���7���X�w�������W�߯'�.����.�#>�_q�\q�q����
F��奯R���l0�J����Ҋ�M&�$��p��&�ż�=}��w������� �=�?�ӻdy��Wy:z�|���ϊ� ��y¥&�_�7wz*�Giyh&I_�6}��h��׈>�!z��1t���<���%��{�H�4��,Ft^��O�SМ�#p�Ԙ�[��*(H��"M�T�{W�:U��K�2?�w��|<b��aE���K�!�L����
�G~1���0qh�X���_X6֛D���u�M��>U� )���[#�H-��0`Ǳ���(|�����]j	�c=���L���B����K�\bm�">�B!(S�h��HLL>�Ma�=�����VƊ�*Ã�^�x�ڕ�&P���MRq�AO*r&#P��k\Yk9�#�>klY�1`��T�����]�?�T���uhHJ�c34� ���u�Cf+ˀH����r_Y  @�� ��IDAT(�(^�K�j	�LU�b,B�l���x0�k)�U����?�.|j��ܐ�Zfs��x�ב�tDhyQc�8|(4U I	��V�!��*TFJ_�Y�n�6�M��۞3�h@ت��*�u�4>C`�4��u��mqm�ڑ#�>(/y�+��� ���.���7���z4'WW�������\�Ul~b��Rˮ"�ƿ=z����Sr����F{�����lkeW�sO�x��u��տ����cK���L�Sો����.ʾ}+��O<�������}�=o���w��l�i!q�7e�;&��;r��ܕ&K�`~�
�[�j��Ag4oD}�rJH!j-Rh�ʍ~�a�%�9A���+LI-�F�y�+!��\�ٗ��3Ȼ�����Z,1�ؙS�*7�
�8gR�g�A	Y�ƱU<���E�q0�Ձ�����U�![.l�Tv��U��8�@�@���$t��*;�#���k��(�ܵ����/k�;�~�t�oe�!�K�&gT5$�2X��4 k32�V�o̺1�nZ���bt��l�X�&���W�`74<K��#�@I4_j��Ƃ�7�d��j��LaP�,�p8�]lt���C�F��*TL-�$�F+�5k��GԂt�2�p���2���8�^��%���1~'����[�̾�2��2׉B2c"1Sgm��	#@�݄bZ�(���0GKjJ&4�3w6|d����"��,аNU�.�q�����Sp��.�A
�31� ���Gu�ǽ� �D�#f�Big�E9W�AinJeň�)��4ӊ
�v�'�<�_�䲣G�����hp���a���X��c��<����M沠��X]�줱�ᨸ敕�Q��o��p����^PC&H)�<`�Q%�}~V0�r���U��_�(�M[�D��m�'��ǳ����d��;��?#_��iY[Y�n�(�de�0��@4��}�ݡ�����Z���bU�L�	1��l]��#Y��h����'v�{�`�1s/`�5uZ3M	�� O��F(B��ƴГQjlc�*R�������[@{�E�Zg֤��[&�u��SH������C��s�1�IoC�ԁ�,�{���P� \Ӊ���ujX2�ȕ�7g9���s��z�;�_<7��M[XfZ��&��|++jv7]ԩ_�P��(V��U�F|0N��g��x�N��t%ue��I�)ljh �ўB.
��#�"�[Ʀ`�$��}�Ȧ�r�֝�XiPT-ʒ�Tt���@�N*j%�������j�f�1+��5�W�M�>��]�1%��x!�N�X3L��2�ɿ4*���`��� �ӛ~�~��_y\mL�	�;vY �P W��ڄ�>\���QT���L�Q�L����tûT��1���7tN`~�Iu����̸�ՋԦ��5cs{�d�9��@�����>T�yy��jY��5C9i�Ңy5毦�N��dY�����~�����-��x�\�&�c�a��^K�lJp��`:W�~��ņ�:�A!l���Ԣ�ϱҁ	A*�X.���i�t�
�>�r\s�}�2G C�n�~��g�)BGRB�N�%2�����-;��P��R0U.;ؕ'�T|xǫ��7�>.��o^I�:n���" ��eDV���u΃=*���	�E�R��dX����a�s=��(G�Q^U?)�b�� ��@K��8���t�Q��\]$f��p@)|X����)N4յ.t����X���j��!���\�l>�>��L����Z��j�'93@@�;�<+ U�4���� �s"ˠ�Ʉ�
���A3Ew2RŮ�WU2�C�΃�RG��C���U�pb��v�15Lt6�2s�@���X)���Z��7n7,�k㸴�/Π����EŘqS�������:�<7_���"��]�ێ�Y���¢h�*|&�,�\d6o)nY��@����=����A��s���'�5U~u6��ӄ!�@�W�W��$�(��e�p�!>��I�*T�FC���==���Ga��6�R2�]�OY�3f�K�gN`�)��l�g��?�A���B5�A��d0,�ځ�ڣiH��}FIժ�V��H���(#��HY_9�@�nvUQԁ�;�Y���il��gjO��b�V���)NNTʔ(lڽ��T�K:��lo�����������6C<|���F���/3[H��z�"`g3������ٮϨ/�²�"[~]5�u7}���7<G>�}Ejs.�K����^�\6��t�Ǩ�C0ne�P�Ώ(�[�����L+�w!B�=C�3�{���%�.1��+�����{!�7('B�[�N�@F3��DFO����i��YT�G6�*�T3U����T��>hs��Xf�l�ه��3���A��B`�&a/_�t�	���m^�!���hc!{�8�	7.a9��Ejjk!�Q�F�c�Am������K�;U��c�-�JY�5
�J�������Ġ?P2�@@�r�̲=(�;�	r�B4��BF�M)�z<��GU�CT�ؘ5���tˌ�HX�+\8��7���~�A%���$Ż	z�����;�"�?�L"��7BR���*��d
ZӏuI�N=*ui��y<W%�S���Ml
W�nn��z9l�4C-���J"
�ǥrd�Z���?u�A?/�c��8eО�3	�j��jo�J.D�1��*��E���`��yE!U3h�|�S��c�[>Xn���B���
���'H�ӏ~�Pm2��Mk0�!�lO�ɂ:�8�4Ŕ�pS%>`G�s��+4Ԁ�Qg2O+��Rk��F�O�/CdZ٪PZcY����%y\v*So��g˷<���Z��syꩋrv}S�����w�%�|t�����G��&8y��;���.��>_��&�I�(�jЙWp�'8��BܿT*�;� &I(�=Q�2`R@�%�-0�5��Fq_�����.�S	�8��-5�fs�������Q���:����6fT��i�f
������G&�̅�.6�{Pp_@.A)����T7^'	�IR���k}d06�|��EA�S�$��ŉ���-�\�oq�7���C��NXa|?�4ӫG^�	9�*?�c`Q�Y��*.6��-'�#�N9�x�^X�Uf��f�)�����i%�"�-�ѵ�<�r�Ɔ����s:٠I#�m���m�Md��9���p�<�`��T�����ͯ����(�	��IMi�e���֘����_L���t��֟1p@������BĨ���m����P�}��+�gD釰/ y�A��fgg��\�r�ml��F���8���'%5�2��A_�(4���V�(��+~�4U���T��Є��X����Y���ZA�RAzQ4w��Sr>����fۥ,��$�䜷 ,��V�-Q�0�	�%$q��A�D{���{��O�W���Q����O:>>��Ž���/N�ᫎ˾�'e�K�^�l��ޙ\}�-�Ol�L�-��t"y�w�@~�7߯�h��%����w��_`f�7*�9���LS<s���-b��� $+�)X�a��PFf:y[�4Ř�O�.����y
RĮ$���=�˛:�9�6|@h�dr�2Xy�D�ڟ�\P`��6�l��.���e��\.�Lt��1Eǘr��d`f���;��c�I�?���!��پ.��,���Dm����I�f�XH���t���h;�=��.�3	e�j;̨�糖Y-P?���E0~���.oj�~7��q�Dݾ�?i���Ա*�|٨�G���4�йf�D�����Z��&0D6��1����Y1�g�F�DR�`~�f.��x:���Z6̜�� ̱t�t�&�*��ʉ!`�W.�)ΰ��f����d�=b�같����1�DO0d۵	�.gc�Xs��,y�E��p X��r�T*F�����,�{̥i�"�G�,ȼ�.0� B���U��xn"V��\&m��G�ѥ*��Y�f
�0����$�T��&�k�F��D0M�,��T�憓�sr�}��{M�cdV��X�߷�`�O����Ҡ�B�|
����B�l^����&�Ȫ��Y��Dj�v��r�t.ם\a�~��o��S�g�7ъԸ'�Y�o{ٚ��R�}�ɾ|�kg�lK��tD4!A��z�Cu�F������l�V ��0m���$�:�p�}�\i�4��������ǼADV�t�'-�p(!do������Ô����-2�PzS���ϬQmH�{���l�$�~Sq�Y�VX�F�]��Pz�ʷfP��F�Rj�ҕ���*d�6�ࢺY�Bn���Qi(�U�6	�`2�J����W�8S�1�O����&�Spf����L��Ϧ6��(�}��ژ�����V����"/�甄F�S.6���Xuf*��>���f#.�m,����+53���l�Dkhy(�%'܃�O�TQ)�j	��4�έ��=�����a�ɩ��v���A/���C�Y%sIc3PD�3Q0s�6,3�q��ѻ���W�'A�T���<䍿�-E��jXc=H�V���z���9<���$�ZL��^�c�2	�=G�	>''*.�oO����� L��`M�JL:��]ae� ��T�\
���3���s�>�&��N���p@wp�J��?
g{
k�_x�>�&��C�׮��U���W^�,7�t\�{�j�@��V6y���_xTN;ƚp	�SĚ[�=��ݿ���ޞ^�cg���5eq��k�\T��<y�"����Ta�;K�ʸ3�	�	��82`��L�Y���3��V�������n��iPk�E��Y��Xe��;6�Ӳ��&�ԁ��9X|i� 'J��
	�)��t�0Ii�_���p��W�ת62.� Ђ�&�5�X�jn_�O��x��
���tu`1��WLAsn�X�d&6�����C��b����TCQP$*v�Tb�4H~��=Rs�qvoIզ
Zwz]u/��vd&����"5�:Üg���X����l�bM�vb:gHQk�iA�*��{�@}O�E����ftaVi�ϰ�����t���TϤ~�6��Ȑ�&+x�u ���5�k�̴S���Ca�2��ܫ}�@�A<��b���=L��.�:{�EAxu1:ͨ��h�kB'.����<����VQIU=hi��@�#($&��
2��g |�(��¾/4�L^B[�2G���lu�`�hm�r��"�~W��z�N�U�ߌ�^y���N���A�H��-�e����cT��A���#���xͿ|��:�,���ڢ�'ŀ��pc].�l��ª��?!�K��F�q��t�1��o�]Ξߔ��+��?!���?0��i���?����0B� �
��Z���Ʉ���I5�p~���/_�Dk���*
�qD�6���M���Wv�1¨2n�o�¦J�mJ���8?�内����x\���sg��e'.�o�oqxgd���b D0�EeT�,�g7e<Ur�9�Fd�a� �V���C>�V��x	.pIK=L�Fu���h&���LK�9YZ&F�LB�dsg��g�;��0jJgk�b�.nKoYF��ZYZ��g7T��Tc����)���2����sЩ� 6�9��p��/Q��ղ���T��\�/C�b�.�n	_W�i���=���	�3����5���L���gQh��g��HW�cS:�?-��u��/K�?��&�U�mPF�0��--MI�Zk�84�E���R$�
��䬣�X!�Ui�x0����8�Ձ�� /�$������p���5��1k`{�
�uc�0:d�aL'L庙j�3�H��~���S�XJ�q���:mmD��)���J���5P��ճ�}�j������a�F���������(�^���Tu��&�ܤ��F|{��9���eג�P,��'���V�,���~�k���d��#�e���s�Ɨ�7�yV�y��4�L�d�41��g��ͺ�k�E�;��hJ������t��(��g̲`�4|�F3��+z]T/�C�$���Svai��®$�}�����h���1�9�+Y
���|@v���=�ݓs�e8�ȕ'�������̇�4�̫I.��7�5d0�z��7LA�	�:�Uf9�x�h@����
��!ۨ�k�����j�B�C��.P,X����K84S�ٌ��E�������������͗�@zU��c�=�,9�3ѷ�ɧ����LO�$刐�"0��d��	��k�:�������.��u�� 	őf��=�s8����_���[�ץg��:U�������h7�́<\�]�xS-h'�nx��YR��ƴ�l���-��p����\%/fi�T���=���S4�yK��m��j4�%HEܑGs�_��1s���|'�cz��{�@)zY����F�u^~?㭑R�|qi���J64����[�/�E�[<M��=���-�-a^�ѳ
�G^�%`�h(�k��Ɂ%�v9O>2��y�{��.�Z���͗s��)K�[����s����3�t�nưb9�߸�D�GV\R��O!����#Sa�dR�I�>kw�ख़��\��)w66؂���b�n�YH�W������X'/�~g�'���O���yû�\Cl8@w��׾����N-�S?���H|���5z��4&++�)�!����ڎ=R@�r�����W�~��z�1V|�ũ��/Z�p	Y!��s7R`�8KM�����v�(��6���VJ����́ ����O��Z�&�{8�*1��E��a�h�z�ׅ��D��0La:��AN�۸��V	��ee�!�Xd���3����{�V����I�a�va³71�����fW����a�LK՜�st�d3TEZb`�Q��DZ��,��3|21"�IDњ�X�W��E
�8��:!0�b� �3������v+�mF��Ǿ}3�8wi�﷚2%����LѮU ���1>9E!��(��̑�r�q�Ҕ�;2W�p���12F*
���f�xk���~�|�����[8�[iL��V�Fِ�sO?oZk�2�O0⛢��qH.���4�3��J�*���h�=���g\$�8�H����4�"f���ࠩ9c�0�U�/�|��#�}�W�&_�IJIT����1�/��~���(g�ʸ�@�h)������&T*܃��m�q�-v7Nr2n����EB(<��3��|�#����Y����JO�x��D��c���5�.E�mT+J����Z��k��3�x����
����p'�:;+���ǰmz��*E�-���Ukg�6/ '�+�c�츃�����˿�*��q�xCa*ܐ�\*��EH�WK$�&�������mF%��8�ЉF���M��ٶg/��A�P��W.j��S@�nj�8��m�EL�d���F^[�ca�����fϜ��I04�������j:D'�T=}m�82^3ۦ���,D4cCuLM*��g�:\F��fi	��b5� �km�_-/�`d�*����C�O�ɝT&�q�<E��gX S��l0�#�<�8e\��i5�`��ȹ'ڨ��c��q�>��`͵��+�̰oÅ�tC�<�m�����-�xn^P4'�<���.[�����+���c-5�ש�u��)Ja���Z���Lf&g����W��tLr����Qt~_���%~�"�����o)W����;D���0IBA�e�-Q���\����b�7n�;oϽ�E����f�͞}̐Egs/��]��q���>�挗��!�2��:(_L:`�i�q�iZ����s���6PEH��Gߋ��U�&������h\�Hd�<c��)�^�%l��Y"(1�FK�T����RT�{71�f$w�p��|c��e�w{�L⸀����O����-2�;(*�V�bmu�6��ٌu1�2�\f��ɒ��pa�k��:.���<��_]��c�)��\��G��F�/^<�������u09Q�'?��4ʌ ��{�y������F,��붕�;�Zgc��tٕ�p����IR �����7>�.|�ӷ�k��&��;�䨦Y�ׁ�
w��~� �X����u�L�_�{`d�/��h��u�z�m��u�����
7<����@��8��t��!��=~���ޅ��)>q���K��%��"�4�ޝS��^���(Fɀ�Z��
J(;YO�澰��-ǎ�*����N]!��3���:%�B��7~�ɋX\YA�	v��?sr����n˯_o�0�"���f(�Z��>���x�N��Oo���s4�t�U8�^C�4/
ֹ|*�Nǟ:�ƹsX8q���y]���aVH�̩�CT@����^VL�p�7��<�x�_N+DI���q���N]I#�Y�9��.��Й�򟃼�Kߛ��$1U��xS�uf�Q�x#NE��/3���+fo�����9$y<���%���#W��u��س.=��x��M�9)�VL�y��p���-X���u����ώ~!����;���}yM� iՌ��E��N��l��-�F{�)6�ǐn�Ȯ�/-�h���Y����^�Jަ������fO�~w��#�:9��������g�;O� ocu>$^Y[�։Xo,��K m�}|�~B~�__q|�X��F �h҄�.S���gW�:Q��~O*2�|��n��^w%����hp��ojŊ�E����!�ᖹ_dޔ"&&�x�˯���9{�<v��􅘞��:�#o}���صc
�_}_��87�Jm"\;M:r�}�p=z�	jd�����4B�v�ϒ����֖U�gtlL����-�	O�
6TڋA�|�m��f#�Z��].���f���Ѫ2[2����.��JQ�P�����+�$I	�B�^#,�a�_���rf�)�����P2[[ar]� :�x�G[:4R�P���zա����Ke�*��RL����mk����L򅋋�q�+^$������˯�d��ё��OЃ�>�S�O�Fq�^v�·@�.|�m{)q� K�#�C[��yI�%Y�5PK�yrؘy��
��m�WDq���#���Q�a�<10X������q[�}�1N�&�s�¥}R��W�КerN�xz�9��j�6�t���#�jXf�P/Os�6��^z͡�j�ǉ�/�5v� L��e�,�N��uӱ�;t�`;�ܽ�W�:;�)�_1��	)��(3���3���+��M��E���R=ی1��s��d��wa�+xVp��{g�hSi�:�༬�3O��������/�Y#���q���������/ߏ��a�5�z��OE�,t��
��o�ݷ�����n���¢_��Tz(s+�
"E���'g�,�B?�K�/>,/�Wjt�E��עȷ:Z!;���B��Ȑ�#��y�sf�ƅ�U������)h���Q��-��oy�!��zY##�C��w>�;� ���֓L01����2�d�0II�A�Vm����U�`m�ڊ6ˏ����\���J�,�H=>S睜��h�Ac�I>*�h�e�9�̉c
ӐI��p�T�%����)6��#w�ɱ�a�IB���X���3ޜ�༝�E��e(�Ș�8��[�ݰs��:m6�Z�������SG�V47�!�y�7��5<��kpj�����~�2\�2�l� ��F�neH�<8G^�U���˜a>���"�L��,���\�Q<6��I���`�,���t!����9��$M��)ux��A�w���L����N�;\i_�"�jh�����Ί�I�r�N|i�3�ɲ���D�c�do��]�#X]A
O�~d�(ol�\j7o��:�Jp���X�Y��m��I�_������5�M���NT�rD�����Q�i�O6�Ɨu��bԴNl:��N�����a9��'�nk袆_��W��>�e��M��^�c���,�k����w��?|?���é3��У���C�$�,v���~!�kq�\���b�y��z�����ݕ6�j���W�R.��#����k�.=���s}r���1����C����0qS�&Z�߱u�6�Cسs+�K���ظ�Rx��Yu�A��rI�~`_���Γ�ރۿ{L�n�� '.t�@��S��ѭ�d����h����",�^�t:����w���#�ș�S�hR_�0��}��xZ����<E|����r�Ƨ����o^�r�����\�a�����h뮪�a��m�簗���߄���!�e��$������r{N�s��˩3�]�g���p4�!/܉��z���۱w��s���\�:���:]U_)*8p�r�:�)ch��s�}��5��ugE�=%W�ݘ	��Y����l�S�������kۦ��Jlö�KA�	���$m�
<�p�g�;o�(x-i���f�����#���Ab�b�ڝ�ӺA��#��IZ�֮â�K$���k=;Ia�.Fw�"2�����������6�H��@��ND8��G��t��0q�R�KZ�%�]7֢G _5=�!g�d#FF�!p������ѐY�IꥧP����4	�C��gxz�g�F��G�2�C�Z�I���>�*\�7��Z�۲U� .��������mxÛ���0���<�	M)�F��٪�T�geXl[�=0cÿY~�+�AϿO�355%�(Ý�.z��]�k*iq�Q]^UǸHN�St�S�m���z�-8;;ON�:�ʂѥ9Lϖ��Y2"=J��!c�u��W�����_��	��=����Xh���.l1o �F#���0�1N;D�ב'P,+I����nM��M&}����D�f�+�j���]m��Í�N5VN\~Ъ	���� I'�s~��L#��J5]`��գ�#qDvi��m�:n^��J|%�Ϸ��k�=R0�WoeA1g�my-Mh�Z:��ԊJwC��-,,�xcn~�cXYY���81-����G!��w�m�_{-Μ����2��D���Ɉ�̞uov��fcSG�9��StE>/�?C�G�T�*)+J���Dp�C%�v��d��{���+��Oh(ǩ���y�t�z��{�=l��I�"c�c�^���2����rt�i�:�g���y�7"�(�ٽ/�3�a��;S�ѾO�z���	��%1H�������4�,��"�
�B�gNz�N~��WS�VN��r�~��OR��x�^���s[_6�
t�gI2���>6�$}��{�u{�..,�YW^��o�=;�cvvSۆ�m�fT�5�����_|Azؖ��4�η�E�!��{Cge�}퍩���Jv�(k���*^{><�nL����y�L$t��#���
�"��4�A��E&�И��u2�s�}��K�����:6��9��p\=�s1O��[Ɓ�����e7߀�=�|���A�QBwu#�q�a�w�f�B�P�쮨����a$݀�P|���t���|��|��J�j9b1�f�urg+KÖ�t�"b]9��ǆ�6��c,s�6�6�Cu��F�#r�]#d�	Iw��Rd��f��4-���YV����j>{ɽf�1�xrڄ�FR<M2�2���F �ˤ�-Ŧ�Zm�
]][K���b?�Ȓ���&hr���d����5�
B�@c<H��u,���q�r�^牷�eK�&���~G���%NL�!�Q45*�=�drhuIk��l�HkF�k��`3�E���P�y����ʅ��e�}3�\@���)���Dq]�����8?��w9.�/gL�@��$���vA'�`�S����b
�y_��{h���9N���vpN�6��n�iސqjF�Ikʛ�����|-pJǥ5�e��_Vlt�Y�x�V�VG�|��\ׯfQ��_}��g�x�M7��o�M�^�>-����mT�>������Y<�W���9�����gj�:��c���ߍ%�ö�����������<vd�]�EjZ#ht�$�����w� �������2>���F���#��5w��(�{�A��q�j�ט7������anr*��{�; i��&�}�7v�M�1�D*
���ve����o}�8uAW��o���������8=�>9"��T���H;��hGU.q�U8m=�\��'�e�Y��
f�j[���B�t��������K(h^/����웕5��t?�+�Ξ1�)��t�VKe1ȭF[�%ۡe�z~�˜h{|la�ջ�^�8�d����-��PY�|t�]�Y1?#s�r��@TY-A�P��*�wN�U	�5]�Y��Bl7q��az�t]C���bd��Q!Ws8%��W���7�-��e�6����~;��>7��E��$QO'���ٴ�]�<qPc3��m�v�a����|�PU�`ɹ�l�C��vW
���z��(�c|u�,��{�f� iޜ_M��
�"\�+f׫)��^���|��7����F�H�ǧO����tCbl���'�d� _��,�T�ű��d��R��#��΂���r,��Y�(٥�<Z����d������nXg�o.�v����'����}����K�{�����/��7p9y��~�{�ů�o����g���s��;(W�����0歠���������u��W+������y�m*��넇�׏�>���}���}ju�w��Bnl��$vo@+|�5x�6����qeA��ey�M�-�0����Q97�1%.׽8�"g�V�ٸf}�&vn���LO��?�_��O��x��(g1�bR?Τ�Ti@�����Xײ�"�n��'iMH䷌�$0^�������B�A6��+�n#ߜ5E��n0�,�4!�(�9�P��C.<D�>z�b��PC4�%&�G�2q��~=��s>�ǽ�-�0�Ag t���|tm,"�4c"�6,	����3��m����N��{�E�wrƍUv�B�X)K���EK~	-t4�>�e��Ǘ��I�ٜqF[̐����lo�^��i�l;�]D|%�w�A}$�+_�-��Q��;�4�vL{�a�]�~�Yr^U��?%��7�߁]���X�ZMc0K�jwƩ�����Д�+~�څ�}7o�q����|��cstR�1���<l�2�$g�b�.��9C�]�}��|?C���F��$���g�]�fd5�Ģ.U��IM�#M�����Q�k���������_>����8t`uZ�����|㶯�ʫ�a��ItZ��z�/ǻ~����F���V�ֵR]�r���2��m�)�8=/���g��o|.=4���	�Ƿb�<r��	Y�6�{x��<��Yt:��^kL�RA5N���ZR}$������Ͽ5��^ c�d�a8��p�hw�Q�=11�'N`ffF��,�G%��>���3����5gE�>d߱�%�"]��D��Y�>�g�j%Q��IX�rNY� �,�d7�٣�4�vh��yTl$�U��9`�
B�EY.q.L�G��>���hbxdX�^��V����)�\kl��s̷w{j��@ޣ�o��� �k����ڂc�Q���T#�*�?wq1+�tq�RQ�j�>V�+�)�x4Ƞlʓ�p3{%�^*A	��󹴍��#UD���Zm�7�Or.m�˥E�_�)U�Z�]�:�y�ZҮH�EH�B��sP�DyW�(H;ȟA���"�W2+/+�9�&��gg-�<l��<m�jO�B�&[��N��%5ej-�t?��Y��큌O��CYCߌ��y��y�?P�\�_��R��|H�Af<��+c�K�e�X1I?�yfFL�O� y�� 0����}cqt3E�<�W�7"*�M�9o�}��3�S!=�uы�+R@�z�2��o>�?����Avmx"����Dc��׾�����������;r[K��=|��_�-��(xb��UT�Ek8>�@���+����������f�!{dhL�4�K�T�^�h����G{�Zh�J�+ۄ�˘�4�Ԏ-��hD� �K^xF�n����"�Ȏ��2}m6[t�iq��~��z�#�<"u)���ݻ��&���=�"�|�.D횢����x");]"�i�i��DQZlo�Uh�;Rhp�/)�I��ƈ��Bj��bEV�4���P`L���3��F�ߑP��B��f;B��۫��W䡇�	K-��;%��mӎ��[�R����m��p4Yhɳ���s��G��j:�77�]!����1�RLYHO���
�*y-Q�^\ZL�z ?6U��8'��*�"�ѬTȳ���W]KB����0-|%�Ş���g��z�JWd��(+�$_�/�cם�H�$dO=w-@ƙ�����sw�y7�ŒK2$�;D�,Q��x��a�9�j��3�s ��H!<�(<k�҉�B�L�C�W�s|JB'�.S����nđá{��٦�(�Ni�L.��C�m}�ݹ6}�v��I�c;C�}R�"�|�䈳<��l�;Y�:��E�kM��,*�s�xY�;-����'c�j���49�:)�W�|�,{,�e�iwt���W��x�;���>��x�k���'g1��*�����K� ����`��~,�ϣ�$Ra��4^�u�'h����'p��q�t�v���K�y�o�����ر�Ǘ�t?vmߊ}�xë��+h�!RA�M^��N�� c�2�9]M�<nyɳ�e�7�J˗*4�L��g=G��&�5d�b#�0k�<a�q�~iiI^[����M�h�n��&Fkc����-�p/��
B�=�
�)&
�e�w�Kck�	��1ǋI�d��-k�1)O1NW���
���+��`��䊸ݕ� �>uۧ�c����t��"G��A����4��rY	�|�"�8�Hv��8nw�����^��/�'���L�hNd����PG9W)e���hKQ�������yLYq��q��x���-^�����s�>��5z��,���wMN�sg�#��x�!l���\Lt-̮�ЙM�>wS*%�t�6�ͼ#i��&���@�	�_�]�%/��\*E�,�눆�\'�I)�r|؛������2ce��?V�8��L�5!����4��+�d��B��1��Cuyb�I��/���Ƨ>�Dyq&R�X=��D�b��;�������|��H�d��Ji�\?�����臋��ʦ��|Ѧս>��G��E$u{�.m����y	�K������O݆��؋17��k�;���a�t�Iٵk'_vH�W:�w�C�=���Wнt0A� �.�q�3�1�U&�k���ߖV�����R����y�����%K���s_l���%�P������O�/S_���^���F��%�-m����񒛯��ŏy�
 ��&�Q
��h��s 9��<m^������r��_3<<,�W�R"�=����|5�����<�AM�k4�W���nvհ�z�x�|8�Zq��l���{Fx���z�&�����������k�u�c�����k:�>C�!�/�a��N`��2�<����DLN�_��L.�e�R�&d[���~^���;�ˉ�}nn;f����׾�X��o�T�X�0{iy]��]�����Ė�4�#�	tSV55آ��`}�"��-��ocǎil�:�ݻ���^���
����<��Z���2^��d�tR{x���9��Lr��������p3f�3����DM��C(o9_�+��rc��v���
'��FP�"��
�0ߟ���ek�� �x�*ߦ]�)Sߦ�{����ߝGI��d('6�w�����8�,��u\��K�'�mV�-8Z��8ʭ��0��j.��\]@�q�ܒt<���sb�+�Ti��y���|m��<���r�x�f�~v��p	�"RQw���F̵CN�?��=��/�W���4��s8wz�~�6��/�z��F���G�˜��\��;b�7A�ɥm���9q�%z=2h�� >|t�ƶ�{���ۧp��2n�v�\��-5���*�\ly8u���(Z�u���w��	�]`1��"]2�4����7ce���*�pG����Ͼj�sA������`#ݴfC>��턖9�6Icמ�c�-�b��=�v�����a1�������Ա�p�cu%��
�f���L=�"�u��DO� @��*֡U��vr�*�V*h�[x���skm�v���X@�HƋ��7��,���t##�L�7�S�b(�L6��R�O�M��=�އC���ۭ.*Ւ�1pn~bl���P��֤��l�����l�+;u�M�m(W���1�Y���'���0��s7,�z�>8p�r RLsK���c�(n����\�Jgb���&3�>�Y�@ޛ�q��M��T�r�+���c�[TK�^�I�_�q#-�j*��;q��Z\��VU�6v��Ԉ��.��*����x���YP5HҎ�<=�;��A��(i���m��)΋���w����9�5u:'Ec�m��p�*�e'��\��d�F��s�d�#Q���(�F�=f���ns)H�t��P��^��h�;��d\?�"s��D����=�!��+Ն�No��G����\v�N|�����/}	��ӿ���/�+�vn��W���������6�JU��.
R�g�"9u�I�z?�y���+��_�O�O�j@^�q���������(�݅9�ڨ�uu|'���~�O��1� �и+|�|�+�đcx�����G�u}l�A�o>E��.*�(T(5����zf���999i��R��޿��?��]h��0^�#���ϦͩSG�V�s�g�s�4�͞��{%�_�k0e�5Q8"ty��m�%Ha�T����4��b�lN��6�5�E�f#$�l7q��Y��s'��T>�_� ����AƵ�JyD�l6l��Fb)���q��ݹ��N¾��sT0�{(�e1��y���8��I�.��12\��*��<��ˌ�cctt�<cz��Dj��βN�������?E�}I��#C��3F[��i���U~ҥ�=�ǟxH�����p躚PR�={33;%�>4T��R�(��J�@}��9�����Q�2k���K��˔�EkѰ����B�u�B�B�τ^�z�v�F�2�a}C�-!�����SnA��pI�H�&��`څ��\q�o��[C��^�=p����qʝ�m���zM�;O=��M�dl���\c��ǳѣ1.䞍B]����7΀ �v�|A4u\�ׯ� ߰�sϡm��$oj6��3cj�@a���!|�����(����;��7���������ц��7�Лq���b����j��goǉ�g�W܀;�C y����3��;�>��\\Ceϕ�y\�b��^�IQD�<�HHº��C����-��&��6N3�]!A��G��CB��O�QVS��=�ْ�����+ќn��~��nBc-�p�l�a9���Dx}�ؘvl�?�E�VL�9 9m%k�"�Q���B��� >��o���	�=�`mu�r�=̝?E;PO]�'�3Uju�}�pc/��d����t��j�Nf�����l2�e�Ĩ�
r$�����E���z4m^:{��6,,]���=�t���M����������D�?1崀n��gλU�(w�Y⨀��%Q�ٷgF�u-�ɐ�@���F�x�Fq���_X6�&*_�{��un��� �v6��9;���81OK��il��}��\�����D}xHr�s�s8D?b�" ��y�5(�6mc��i��3·�F�$�%���<�f��{Y7_������A�gѤE�R�n�'�צ{�L��hln� �����tIj\}�X�d�:�����ޟ��oZ���u�����E_�a'i�"cN�
�A�o��������~%Bu�AX=�Ƅd�X9��M6�5�W���rK�"�޶}��G:A�T�G�1M��Vn(3�5�y���j���
��aY+U�N���Wh�:42�ze�wӿ���Z+���>��{��C��K��u����GN�Єp���˭ �eMk��=A#m���}Kŕǥv4m�&�D�BC�n��Y��*40�W�4��������ϼ�e�iп�&��|!���"^7����*ǘ�U���?s�r��k���K�@��� �^���7r�HPd v�܅���L�A����M�nSO(�<�1^��RLt�����r���z2�|)P�m����ao�k�l�_m�<tȀ�w+t�d�&�L�C��ѥ��\�	���э�Ŕ_Bb�X��}�^�'S�T��I~mbb���-c���Dϱ$*(kt[*5T�����9ɻh�$
h3��H7T���:F�������.�v�>��Z��_7��������_(���Fq��=Tj���)ꁄ�4!z*d�
�W۳|����Ԇ�՝�C�9(���z��pm+E 8VA7!�X�-�ݸ+VȢ"��8|foۅ�B}��	��"�_U�Ҽ�m���⦐'9�TZ�a����J�dG�{M�7�<6�	HGI���]�vb߱�V�� �НוQ%��_��,�����r~jT�����bG��������=/?Ɍ�=N!9�k�!^���֟����]�Hj����ǆ%O4��d\Ն�-X���7��;�ex����~N�P�c��;y�q:p�DO��G_�h	..���F|�+���4���yTˊ�`P;l$�՚��)`�|��dm]rpV�)$�c��NW�B�z����cH�4�"��Qv�.�k/ݍ�~����~��xĠ�3N�wE_֗�r�h��.�Ax]��	�Vk� �B;�l�9u{�m�_o;O�~+Bޑx���M�:yW��{�~�(�ڳc����'�� 5|�hGrۊ��f<W񅔾����qi1�2��{�]�q�8���e��0@�M��JM���}��ٓfAN���F�HW�3�(0=]�+-Lm��NB��=_T���p3�R�o��A��=2�Ò����zS \�l��<ͰI�~?W��r��b	K�k���;kA�C(��bf@~pk�˯��/QV�,&4�v��{dd��yQR3|�=xH���?.��.��cQ�.zZ�s�y����`4����Y��%��v�Ҵ�%�R��@w۬�/�� 0Q�L1�Ǫ%<��`R$�j6����<�ͳ��8���v�I�"����ƧE43�v�O7��ىG�wj��NN�ɍgڍ��b�o��F����}�3�%㔒�[On<D��[�=�b�pmo���\�?�"X�|{�R�$ �����U�ƣ�U�bʻ�s�ǣ d�\ԇk"b�R}E��j5�o�~W]�E�-8u��К>����	l�;}%!��}���5|�wI[��s4.)\�&%�/T*j���bL��E����r���kE�>�1wy�JU�%b˃}v+����ѡ�d.���tVgq���E7]������*7�~	#FD�����RC
�Bpdvn�s?���޺�����&Sr5����Ù���. �L"���aS8����8~�)��L�=v��OiVW���Jf�2*�5�}=md�7�*�6���)���H���uA��{��N�����rYQ����S;D���J�*^+�=9���*3@�cb�4�'�G��+�.�f�n���I���$�J�"y�c���S�qsOQ��"�ʩz��T�P�;��:y�m'�B�}��g���Vuz�����A_!�ͱ1cA�Н;�`�B˵�(XK�5�Ǥem٬�(�����i��b�m�9� oc�3ʥQܲWh���b��p]S��1����*�)4n,��̄���v}��2)�F�3���cA�YC��$Kץ)����H�f�74 �O��2�iK���2%��d��t`7x���l6��� %pj�`�o�Y�vo}/{o	*�{i��
d�~k�;��y�Z.d�xg�Ew�z�
s�5#��y��;S����ubHU�(��w����1"~�_���.�YƋ_�l���O<��)���q�C9��~����]>G������ޔy�6����~�Fa��q��&F�1�Q�5���<��n��Hn�jРy�S`u�O�nUz2�;��XY��������撧�F�{8�M;���5���:X`�gE�6����d��Z��	L�E�j�'F|4�V##����Ea��X[[���E��d<�4���tc�郚�U�U��;�
���s� ���ubt���G�H�P���FIȃ�ŝp��D	��+;�jc��@��a�mN7��q�6ې�q�0�N�Z|Y�����gǆ��8ǆ�q�R����n�`�(>�1��Y"�Z�h���^E�ZQK�2y�k���t~֊Zu�\O A�p�A�j4Ȑ7�@���y�W�"���bv#�F��
s�0�d1���Ƀ���J�#��b.�H���#�aL�o�<�e9�!�ƒ��H�2]Î����K˿ҥF�����"!�4mQ�%�=�����["���aW�%�ܾC3p��R��D1l�����B��y�J�Ǡ�)�k���������tX�c����H
GU�`���͇�-�W(׼��i���V?H��Zy\cL��A��yܩ�v�0��$+n������I9M�����Q(� �P)x��H�Ӎ<��w��D���z��}Ë�o�+v�b%�'p���q���ލ�F����ɓg�(�0s�ƨ�V�o�����Ǽ>Q�l�z�l������l�?�_�����q��9�����r�=��s��
y�B��@�Be���@F����f�y��1=S��r��`�N.ۓ�0�������C�Z먏S ϗ�)Q(0$ '�����r��V8����������kɫ,*D��p8��ڢP�j,ˉK(���YnN�<{Ѽ���ot�����8��\������I}qqYd�lJ+��;n֡�Gn��|M�0�>,xR���4TD�F�lqI�z�I8I�����Y���h���LQ�_Hs�6@���°����bX�R��@�Y�ȚBR泾l(<�_�r����(���Cր�]�ai�6�y��� �p���d�?��ku�S��2$�;/͞�y�I�Sȡ�P���4�#�)E���'�Aʝ�g(���z�=�VՓ4��6�]s�������g��Tb�w�$eY{����sbU����1ƺ�<��ޔ���k�X�#�2o4�-��@x٘���.�{�E%� ]�bč�f��G�ή&�pg7F��[qR���7y)j�~�sbc��N�dd�\id�gR-W��9Y?z����AG�T��z�̐a���!|��{���Q�M��|n������ރƪF��O�E��,{��;�E��u��[y��°�[w-�n9��߂�'/�Ͻ�Ǫ�(��~���2�CG��+�q�����w�_�G�x�����s#j�&Y�M�k����/�>�&��S�{d3u��;C\#goyM<V��5����p�GkP,p������a��B�8�9O�]ġ}�ؿo+�=�U����f�c��r]�pl|�G���V�2m+Ϗӑ��f]4_��^�T^�����c>��E4Pz���a�7�O-3��,�ki��FK��J�F�[����3����z0.�B:�E��'��1nWw�w�厺͊S7���F����
%���dH{��s90�a޵1(	U��X+P�&����e=KȦ�4�C&����_�DŚ�M�P�1Λ~�e����%I�ui�:6lw��=�S�9�)MF�Bɞ�}�{`p�Y�3��Ѯ|�z��(��Z�;���;�ҩ�^���0g��NS<s1�9�Km�M�z�qJ�
�[,�����>w�<���6F#�?nې���K7�8�؞�|����yf9�]~n\�ሣ?PN$V8���rl�l/Es�V<tų��i�� �1��?I7�$-���X���,.��œT;+̗��=ngw��G�|�ݔ�c�X?��oH����O;�ŅvL�k'�{�~���?���V<q��@Q�6�E�F�YH$qV\����WV�w7{�c���~���wb�.sz�x
1"�yÕ�`�<���ý�>������������m��M�h>MN(�
�9u~�^?�sg�s�~�>��Ȱ�����쑱W{�oq���T���ЈW�)~`M���"��_�=2�����:�56�J�_\�7%ʉp�K��"��H<��.��Z���PRF�EV��P_���0���p�/Tx���E�����Ov.S�x�e�=�à��ɠJ��Ј,mA�1<��)�B�p-���)�^>,T(��;,���kI���+ya��-2��~Ӧs�(��� �6��2��م��'t�l�����!���"E�2�n�A�Q���@!VF����XoI:�X)clbDQ������:<�TO�9%��)$D��N#s�v�i����G�9�O�#��獵g�)b�I7�i��3�ō�+�i��c`��r��P3���l����6;��UdcJ��Yr�w�{d;��M�h%��l4���0�UF<���Ԛ���Ɔڄ�.���Lq&��R�2���j{���h�)��q���'��&�	Rp�U�����l]���A�[���D7gv��\�!��i�Rs�g�k��V���$/B�$��d(_���������~ۧ�ᡇUf�/~>�;�s�פ	%��� `Gi��p/{�������_�\���j➫'�KKr�a2➧���3��.�B����&��57��>�<��QT�3h�<A�pm�A��î�g����x���[
c���[��xNN���nK��X]:�}�j�ɱ$S�k���U��}�<���x���Gn��*9��p;���X%�-�,>$L��S��5�;�����yr	}e�����a�����b �I8�g��ӉQ	ɰ�"�$��&�{�6"gE+�B	�Zv1�u}��"������Z/����b�/0����Blx���H�`UJ��e/�ݑ���A�6�0��q�Dd��"6c�K�;A�B���C=�p�ЧW�3�q���u2�=A��e�&��1oJ�6��=Ԭu�K䍩�#U�4)|�w��������d�]��3���%) R`�c�h��a��w����F��/�E[��'�D�[מ�I��6q޻�i�h�N6�3���c�s��*���70�ω�`g�TC�{��{�/r��h���r���'w�3v"o;��MMYJK�3���z]ÎMg$)dR�;��ܳ�H���{�9�=�4cN`سt�[�ۺZ%9'�]�����[��N|�Qo����K_�&���+d~����]z�Zr2��a�^�ۙ�=�~�Gq�<p�7�4l��5T���&܊���<��~�5�(�S���*A�ss��^X�ãW?��(՝~����'fq�n��B�Vfs���غ��Zo�zx�'�}w����[�b'N?�8�I"�*�z�s�I?3d�وQ��@��z����L�w�s�I�~�U)
*����9�)�hD:��z>��b_�5�p�4��h�bm�;[n-��E�<�8}�lx�J`R>�K�mޤ�u���Ī��Y�	|4�&������E1����R��0ᜧ�p���K�k�+t�����l���6��6�cO'm�Z̙K�=]y?+_$-l+H���E[]~H`��OJ�4*��vEC�E!��#���+�[�djR�Z뫨��I3�<DZ ����<�,ܮ�e?JS�\���Z�K�=1�=����s��D�u=���M���Ā�'�B�gg����m���p�����HZq�XXȯ7�f�����0;硤����lG8�eoՅ��<���������
u�إ�C8�SՑ�� �qҸ�:G�%�=��C),��v�����fQ:6۠C�iӰȵ��%A��(���N�v���^�@��5�\,�b��$9;is}�G^�V�`��`چ:�&ˌ��%l�9���̙���m��9�{=>��O�����GgE�;7�pD�xǫ1�c#l�㞬ߐ�ѣ~O��]{��������?�8��q�����v.�=�*�!K�dli=r�s��1_���ict���&.=���� u�;c�fT��Z%����1I{������ِٓ���8��9l|��#XX��Yt�1Zc
�Hlc�WQ��rz ����[�om�me
�z�g�^t��6��ȸu����C�Ͻa/�_\ũ3K���2T��Ը|��Z+��b�"���@
��_C1�u���vy�%QҶ��^JE;r޺�lK��;����=�y(�D�o�Ɔ�ղO�7E"��`�'�#�5ӭ^�։!?���i�h��)������?���XA]�'JCD:}��Z~���, {�h�/\E�z�*)�& ��<r&�q|��Wj���9�n�N�0��#3�.�$�f�^�aO0�R���F�8ȟ�X���Y�`��J;�t�f�40�C���g�#���nV��(��=����\�ۥ�)�ȧFla�I橋����Ȑy/;��Qm�3�"Y�{�ԛWc�4�K�ن��^?s�a�3該N��Z�/��H�V�α0�5Rm3w�YJDܗ���fexmyƑ6ܨ>�^��G`����������Xx��Jv������'i>6���#\s�>��[���� xX=X�G����®��>�Q�͐���䬰���˛IJ������I�{nvw.`nN�����p��Qig����YS�=x?.9t��-X?�W��CG���Z��.�D�ZǠ�B�f{;��S�k>M7~A�\�A��<����r�ȁ�ئ�M�ژ�^��S�pq��۾}?V�)R� �d0u.���y\�g��S�Hd�`��T�J��}p9(���Z�BIg�p�>�RJ��b�^W����o�{&��q%B�<ξ��o�\�PԍW�G0r5�blW�U��#5p~*���"�y�2,��D���j�y���&�B�d%XXma���$�R��3� ��u�����<.�?����o��p�V)l�`���7�1{a3ӣ8vr��G9�ª���Uk��R�N�Q_)wcу<w�I�G�p�y_ffd�I����0D�d�����ڱ�e�]f���J��Z�81�%��G�B������Sk?�߳���3\���]����~g%5$�L�Ċ���"(�᧿wi��������~���87F�>����(IR�S�6˟7M�gQΓ�P9��6K
�=+'�����9�J!�:�
�&�����RFh��D ���<�|��	���i�G�����Y+z��z��<&q�b/�pjA[e <D�!�Bkʿ���#�,�_���>�'�4Ȱ���{=2F�}훸�����*�h~���#�;Tba[�Z-��F^#m\u�>��ȸ�R�bO������B�}�n���=M��v:W󋋸x����t\fO�Doq~me�1�;Gh�I-���*�цD��h����ls����RG>��ݳ�e�WOP`|�i�{�Q�{��x��:��n��k�9VGP����>&'ã��m�0u.֙�s��
]2,��2��>�������T&��.�Q���
�χ�k��z d�p�-z��
�����pwi ,��9X�-E�<F�(e��;C���� L�u��b��m-����'��q���� �*<N���)� J�>��&n[F��A�юp�;)zX���w�dЛسc�I�3���<��ۆ1���ѧ{�4�}��[�W�F�q��i�=7��(Y<a���p-���Ϛ�/�@��&��}�~�!�-zs��t
��C�?�g>s��������_䫐㐎d��'ޜ��Q�p٘�So�j	R�K�Q)`�I�;)�g:X��:����Aj =�zʇ�J�y٘�{뒗,�q��p�8��d�s���I�^�����$_xi�%��b9Xb���KG�SA����W.�ȿ��N�r�BӜX*-��Ytk�7��9�n��0�q���령�@F��'�<M�� �?q�y���E/%#������k��J��W?�?>�_����?�y|�Ǳ>�4V|�e�p�n���/���)��r�`mI�-�Q���><"�O<
[�m��3S ���H�A�o�ޅE�G-�^<��_!�S�<���6V4ϚN_���/�.���Ӌ1����}�'̎���ԙz�C��=ۦ��{,^4©��@��3b���lB�>�{�v�BR�0��.�#Ȼ��0�!0�~W:�.=���1\s���j�������j	�1.=<M��}���8�o�;S(2nX?��#�`���i�R�?�:
�b�aS�mR8��f0���<-�*���v���HAȸH\�7I2�-M[��rB^NƻR/�x�s	���yݲ8/_���j�i������O�Hi�b;���XZ���.�9�S%�=�+��
q�A�p��:y���3�<֣��Wp��i�R��n5PV�Qw󙨰{�{G�M��ɻ%y�NX�̖��F�][�!+<5,�X����a;=ظDH�'�9v�յ�ʧ{�x����O5i.y�9+����s�s��ޑ��Iv8������"�ըGQv��߈T�Y#<?qc����A�"StqUv�j|sŗ�3>����Lϗ�ݹ2p�z��G?-��5�wYjE�?�H����S�d%��(��j���I�E�&��x�H7m�pMf����B�\fHgv��_}�����{-���{� a��u<��<��Nm�����>z��]�5P�Nbz���:�;��5��IPg�GЭ Xi�f�EQ�_�F3��-�r�)T����o�4�{��ՏM��LKɥZ���UNi�kc��a]p�d�1���^����$˙f��Ǆި��Z�d������3g(z��
K���d�c3r��698��k���al3�J�"RE���rN;�@��]����8s���;+x��Dq������W`a9�̖�2F�����YG�[�P���,�yj��2�{f4��?��u֡��m����U�=�����X&P�\���yp��V�W8]��ȓ�N�̼w����?.MB9����0V�����LC��J�&{(0���r��,����=[qvv�v�5,�G��f8n�ٗMai�)��[)|�I��;O&Bmx;=�nZ������n[�~34��[�X�l���������#���	SP��b!k���'���_6��1x7��p�{�7�33�#M=V"-i��;��tg�ic�D4Y��&�#�8���B.����n����ץ)"'z��=aƌs���TuFSp��s��v���b���D�ܹ��7���Q�n9�p���׻�[u�3R��	M�D35�PK_�W�0�u��b��y	m��WvON��p�׼Ipm�7���k����G�k*#[�F^���.�[�zN���51]ǅ���K.��;������u;5�}�߃���?F%pny ��#�-/�	N���h���+C����<�ȩVZ{e�z�1�#�BU��>�����Q*k��*)Ŧ�J+��X�Pw�B�o�sS#C8t@S-��q�Q�&�6:1N�5@�cnnE�~��,>�;q�p�w�B�u��#)�a��	��6�;~�p2��@)6�'��jъ#��v-d�^I��]����][��~!V���M5v�ҍP��Ѣ�(,+$�6h��w�.������O�W�(\�n�8vӿ������]
I�.�HwLNW�L���2�~L�͘⸟�x9����f�0v�ʛ8R�
�������4�Ƈt1���Z�Hc3�<W�ȣ>��m���ۻ{�E�s�2έ��ܢ�/�ֱ��)��سc[G����w��:�J]SE\�<w����&�/�Q�AƳ><�6��͵��w�B��4��b�*K����LŨ�Msa�ll��d�޸�
)7�&�Qr��a�&"�Y�C�k(�t)�ኊ��\�.Z�I���5�)w��ьw��C���w�)�8�u\2�%7*^e����N�2��9��=�k�\T�ɵ�Rbè
R�~p�gL�z��{x̂�j�n�\eh�m�K���{bu�lx���T�G#�z��� �[6"L��!��,�L[ B��'����lw���K��7�O�Y�9������_�?~��ƙssx��~��'����4��Ɠ����/܃ �@k����@��j�Gw�#y~��/���41�*4�.b��BZ�e�g.$����Z������{p��O��+�1��'��a��g���CHB�uAS@
��^ji����kx�MW���9�w��^x�M��}�����ftw}�������=�>��bѡk���LX��"4'�� �Z9��1�!y�R�p�$7���ڸ�����ۂ��|y^l	11J;[�<.�J9�8����Ȗq����¶)M��F�qgϯˎ25QC��m���׀m��^l�����!ꅪ:#w-�Ī��詡�4�@ȝ�TJ���2�4�
�Q�n�<[������q�Uq�
y���<!��E���4ʵ��/�y�6N!�N=A�$9��Rc��I�67�Uϐ�>;��z�eAz?��۵Mg���<#Tz� i#�ɵYϑacQ�u���3���ƶu}��m��N!�d���8���E���og� +:H[��qa�c�cK˹���0Ȫ�n��?5�P��[���\���>O�� ��51����\V����.K�)��%N����[F3�]"}^�>Z����?'��Ȕ��H/-�:�_ddQ̇$���8^AY�j�e2TmC��JuEb�6 ����6�lh�����DI����a�h �$䡏Ol��=�������=_�����7����������-��C�;�n��m��2 [�*��'�:d�0@�W�Ok�ǖ�K?�|x�+�h6v�����7:n��J���ƚm��U��(WkXe�xCqW�s�Ǫ\�"��(q}�TT1�,9���~Y�t�4��G����3�0��f�Ա���_���=t�P�(��
;h���H����*=/%� Hm��H�)t���:t�%O۰WC��W����N��r?���� ���w���s?�����煅Y�fg7��U�Jm�.,k��ފSg���pyT�W_�W:o�w�^�,�5Ĭ?�d���*�՝j�Nh.�F4l�Y�F�\'�@ֵ�Rh	,`�-�lO�x�wu��E1ܣCe�h;�4��nI�8#y�U��%��M�"'Jhs`i����^�{t[=��
���+OMI,\qh�_XV��U��X�PgL�ؠ2$��	��hb��d�I��H�kW؂M�ś�g�3�� f�C�#ȸ�A���]�,H���S�I�ڢ$}]�Ph�O�]�"��FC;1�j��X��N��i�,yCm�>�"��AHR�X�Z�[�m%~�Hq����|�׎Q�9�������wu��(��p^��#����=Zpu7����
�S��`�B����i���[�E0�TM��9�'��iv枋Ԓ�"9`Kq%qEUh��m%n�$��yu��v�~n������ގa��O�����Y\y�%��?�k�۩3��ɿ�á�7���|��Sǁ���/b��
<rj��F���=�B���/�����͐�����S�b���r].���)��Q��xxD���UrV˜�n�CV��m�#~��@r��(͇���=�u?uN��٥��9�]�b5<��1�-u�ζ3,��)��f�z�eEO%T
U!�b�������m���2ڱ㟠>)���ō���q�&�֙�z�x�+�Ƶ���P�;�V%<iwi��	,������m�Es��W߀�����z��T���p�Ǒ�OQ8@�#y��S�t߽{7�:y�^C��eL�6I��x�E��,��pA��|Q��wa |	�r����A[[��}��ՠ���N�y����s��n~�,v��^�Q#S#8�]���z/{�Kq��o'{s�U\}��`��݋��7\M������P�W\��p ��,.Q*-d�,��nY�l�"_����(��'��7�u�+�=S3H�	ԍ�%9���'�P<La�o�����4#�h�� s`^��^�Kl��9�Uf�6\���[�Y�����%=�][g��)/���s�)����K�#6�;Ky9<��v��kө�yXlD��o���r`�6� �>�q�*��9a�Q
s(�I\7�/���m��"���/��.ܞE�S��@x��9�T���!oT^�*��@E� �5~�``]�^.�(�_�/c (4u��&&�+��'��?�U���ށ��;�E��^w9>�?�����\y�6�N�~�^������qܭ�̟S&/~����Ƈu1Z�!�"�E�F6gNӅN�&u�>E��\2�0SF�����][OD��W�0���N�")%fY2��5sM��9����Ek��Dd��� ��h	x�	�UU�+j�y�%2�%tzma,3���H������^eM_k�N|�bc��5�♔
��_��O6�{��\�oC#\�h����À��~�#��dM�4�:;��|�sx���l��2�oÉ'p��1LLϠq�$������EL��qf�Iռ��<ʮ!Χ9�P�N��J].W�Xo��/��b.'��*V��P�^��<�u��G�{��qV��gf�޶�jW]V�,7l���1	�B�� �����~�@I.B�B ���T��\dY���J���~����<��̬��Z�Wf��=�)�y���=o����I�.�id��m��<]u�3hσ����~rm�v=��C�k�vj.W�>�����B���ɣ�i�Et�����k���׏��Nӆu�򠎟^���8���Q�����q\\i�5��fB�nF%f���cOc���^Ul4�]�9�oF~�i�w�|���`ߍ�L�������R��#YP$3UC�[���	��c��e6,�`�x;���Q���V8�O��%m~�5)�Vu#&�K�־#0;~B�d�� �^#n;w�9�&Nke�s�b�Oӱ�!�J�E�^L�I}?0�X�?MG�(�lW����Hj�^�z�V�Oi� 0�gO����|�o���%�Q 
�9Gq�mvL؋첱��d���0�~�Ȧv�UW�7n�����>@[�m�?���	
fS\�я��q���9��ՒmcCG�ѯ�ʳ	0j�)�����Y�Q��B�ɘ�f���C�"� 0� G����'��-�U�(�*���B ؂]a����>e����(���;j�T��F�fQ�.����I�'���+r���:MŁ�p)t��Rl�Ԛ�޵�6k�9-,��O��e�[��L�O���/&��|W��C�(��ч���1��e���cG4Ѿ4_���N�%�w�歛E㰱�L�z��7�:�A��k.����H�hz�'W���2�["�u��h(t9�Ș5�5�5����F�X��xL�NĀb&J�:����c���T����-���lj�|���'�<*��v���s>v�(-,�h��xz4?��v�|�ʹ灟Ӎ/��,������_��|`�A}�/��-�6G.��o�k��n�b�x1~�)�������Ϣ��I[���_ē����չrE��C&:pb�����m2O�|7a��<nďO��7��j��Ƙ(�7�Q�T{�M�,�ɝ�V��XӃא�L�&�K�
o��G�
�N"��^h4$-��� m�T�w*]��_/�Z#�_��<�c�0/��煚�1�����K9�賒#7������G���y�Rsb��@d��i�o�b���u��tZ��L}4��P�Y1���
�cK�b�.��ǾK�����:��3W>�b�X'�a�w}� ��;�C�_����{�1���k�����|�����ھ�B�Q����;B`�@�Al�K�����8rx�n���t�?���tz�=؄�=����)37���x�����W��^h_H���X.���ؔ��B��ҍ����H��O/��������b�����~����>�8�����W�/S�S�����t��.�A#H!�tD�w�߼O�妲� ՠ�[v���� @�!5�Ӛ5St��?&��*����J�N��كt��a�������_�ޠ��������1��}X�n��5�>��x�2���h[
�)a�,[�к�����NF�C�y�h���g��d���>J��$���Cn5����5��t��6�-�5���>��S����N����� �t��1z�^���q��.�/���o/����)j�Ɓ�5�x�S�J�K����j\Dz!��J���7KɣDޘVO�<��h >�mv314o�WKQ�BRV���:���_ �{��<�}:4�Aڤ+|��Lw7�D��w�)�F�n[`������9��O=p��"=� XR�躚׶(xs�*H��C��އ6�h.ۖS=I��ckG�4�ؑ@�  i�Έo�S"7i1g㒎�ҫ�����XT��	;��.;��D�钘���g�U�`	n�6B������!�r��|C�z�zt�Y��߾I���-��>|�oi6�{����
@ T�ɩb$�[*(�v�ϓ.Q�\�{~�0�?v�^p�5t�L�6l(�A�I�?&�w�{)�i��>ur����>ڰ~�������NY�K�u���Kɤ�4^�F��Ѯ5�ͱ7�;Ԯ�L��'p�=E�v���Ի��R*�-��2��q�\"�y֚Ք%���>&����Γ.qX��ѥM�����Kx��u��|		�LA);l�Z��>;O#�t��))�߿����������ݗ�OVVV$��R���Hk�����C4�a?s���j�s}��#�9^���Z�I|G�� @0=�dS&�"J�\��Fߣ&vlj�� ���z�3w��X�z��W�� PB����L�2G���c6��\a��~�nZ79*�dzf���M�eD���Gh���4:��tk����in�A���5c%:v�CYx���`t�Hs�e�265L~w�29eX�"�؂����(T�f!.L|8�{"Eu׍����X� 6��\�v�8�����iEr��3k�X�)4h�h!��,6�9!�R�j:����
ۑh;8����T���qvڌ��ǂ�]���������lb]SxD6�/�ԇ��gR�6s�#ݑ��h�
D�suD%���i�
2I�_!�9Iwb�=7�$�M��n٬1�(b���q��!�?C��^M�Yc^(F�g�KT &ßn�1�7���dL����x�U*���u��0���/�o~�>�ܥ��ޣ+yv�-��E����|N<�n\=9j�]B��������"�Y\ p�tzm���+�Z��UW�z�ha�G��~wm�y���S	��㮻~FS�y:~r���{��`/�Gi1�}�5�Lh"Mq �:	f�%lhW�-��,�s��� �'ъ#��8���>�,��{�x,�3	�D.��.���PY}������r�}JC ��l݄~ѻ��<�2ۮ��]�S������CЌ��Ą�~��G�rt~�ʆ'���f~a����q�f���ozc4=����R��B[�O���$]���Dt@%�z�33�TםU�I�"�+��4�`� 1L)��A�"�Z;@�׍���y�~�p�@r��0|�x�_�b���]�sO�β�}��	�V�҉�)Th�ŗG�P�$9��;w�����q�vҡ�'���x����R�̛D�S�1��WFH�l��lJ�T_)��D`����qY����]e�#'�$��- 
V�Q`�� �Y�x�e7Q0��}5.�F|$�<0j�K���\�W���4*��F}"Ԃ�ܟ/����\4r���܀��4��M����r��mpnriQ������p$��3��eA�R_�'�B�Үo�����!iS����d4{�{ؕ׵�G �(\�x��|`a|�<��i�o���kְ�A�/ٝ
�
(Dn�������$V�:F��:��w��1@@��4�HK��%����c��ަ�\��p�OS���|�|n�<{��Z�.К�1ʖ�4���ޫB��)�p��:�}E�9��Ώ<%�٪�I��G���s�u�}����D�wϾ3�s���=��
;Y+O��<PEҺD�#�%6�@�T�s���`�D�-�13��XH�V_�'�"��5BEI�*��l�j��ANipe��B���O���E���>O����yOyk5Zb��ԩ���gmҹ����*�)��Y�А�r-щS�����u��I�M[1�`\���2�
}��K��Mϻ�w�"k f*S��.�A߸�Qt�B���`B5_����Qȱ�D�V�3�_&�N�����eC@�#i��E�,��l�@�^����i%�r��ϣ�ب�p��\�$�VW��f:l���=�YZ��r�"���rɑ���}t�䴈K���\��y2X4x@]2yK��#��i"��	Enm?��☝!jԞJ�.� z�1�a\xSNlǬPwu����O��8����)%��#��bd�m�I�	~��F*ڄb�;i� p��t��5�a�g��ѽtH°�Q�!)6�+Qc�E1EOx��_�׉S"�yT�:���"�!�暄ZX4/5��i��Kcc[��R���t�7��4߮ۦ5���� u�k��6����٫�����E�G����<3����eI�8�C�A[���1�sE�D��@l����~Cg����x͸9h����U��ӆh/'Z�q=�,7��42�N6�BI�+�h@���&��z0��"�Ӓ�ni�MՖG��/���\z�>�|��v?y�u����4�B�׽��TV��T�:�mK��`�D �L�n��JW���!,$
���S�l��,!ݒ�H,'��]S�p�߲�PO:a��|W��x�)v˾�[����t�'��ѹ���g�Y�[n�P%W��O���.�y&hq�SsR~������st�3�A�x�a:��64��$E�r>O����~��t�+_)����n���8��hM�K��m	�d�a�8d�lHh�m2v�c&���[H��F�t:����������Uz!�+	�Ps�>]��+�?�x�GGy��ә�'u<\��C-Y=����D׿i�&������iۖ5�}�ͷE#�/������ѹ�.���5
9
V�y"��$����ѡ�����%���N93�Y*�=�a�����Zc���0��������P����}O@bJF58�>	��^p�b��@�⤄V�J#-f��z����M/Z�Ma0%av7�(���N1��Il4R��� ԅ�'2�OxF��q@��hѲ�g�So#��t��!�4vQD�$��B��C33��,��,Οqxj#�z�|��
d��X2^��JM� �>99��v�ж���ܐ 2������girjH�Z>���:6� )���ma2���������#�#�5�GO��$\�b�����	������@��2�P77�r���1�&��O!�@]�*-��5P.Q����ƣ�H����<{���8#�W�2GM>0s=d��L�^�1p,��/�n�X*�S��ϸ�UNWp���{�� ��Fw9�W�6fy�m��m�]H��K����u�bL�
�#�F��7(	zx�9�rw���y:�I_D�v|-�Y6
!M��6�])�e���4w�,]s����/}��y����-��r�֡e@y�Z��.���$��g?��g�'�8�a���Mq�D������Ӌ�&zr��R�s,�E�����\�-��������U6?�8,�N��K�~��7�Cn���	���f_8J:p�FF��877GK��?6@�3[��ӣgs���#���-������F���$-�a�~�g�hl�L'�c�ec��h'��	��E��
NW��/�-��� �h�U5d���X���T�FaJh�p�'�|�7-�[s~��MSl�c/[�F�܄�J>:��`ۜ��5H�0"��Ok�1$ɋ�/�;Lإ9p� D�n;�=Z�{`s�q��yQ����C *�ieldc��Ƙ�N��4~�0�jc�g�^����S�x����l�~��OiblXx���~і2ϫժ�٧R^o(ʧh``�Μ9#�3��(�%��T�	Q�cZ���>3;Kv��W��Qq1C%6V�*Q|C���KM�MX2�@8vsM���F��yFu_6�(��zYJ���y�$_Ka�"�&H?��g8�@P6�
ziTl�E� ��؎瞬S�@E�
��~[V����!�Yne6������O�<�|g}W�N�Sz���k*�Þ�`��bP3ڳ���~K�#CnAm��2��DM��Λ��F;5)PByf�k"\�2%f2y3�B�e���р��h�QN�ˤ�`g0(�E~!�rf�FJcl�����Jw�O�n��!�˞�(�}���K�R�������+��@��m����w)*���y�x�vj�`�3l�|���.��;t�ܜ�u��
{��b|���BO�	e��/�BN��
�'��9�I�Ёf�o
x�\@����hlL(����wQ�������6۫�p\�?M�J��՚��48>���;.���������8z�M�k
h���5[���:m\�б�%97�.�׆��op!�rQ��p){&!,Gx��nSQ��!8�r����6�b��j5�Yo��h�*��zC"�|�y�^4TΏd>[�K��j���(�x�J�cP�/pL�z�&-$�cx:�˲.^ur��MŨ��T�p����x6�M_p"��ș�DA����k_�T���Qڰa-/�z�HMʵ��¸v遇i��6�=Q|ٴq-�� ]v��A:�u=_r�v3�&r��c�_;%�S�蛺Ț�	:t�5:M*��蟣;6Ja,���dP�IJ�]��C�Љ=xרwK�\_��РKT�5'Ij
EXuU U��Xd݂*���5�ꔬ� :S��أ�Y9������n�>u���(�s#l������+6�	��u{����Q]'J�ق�cӁ�k�0N��I��A��k�@;�16ެ�
E*�]�����r���y�d��c� ����f�k�3�<�]���Y�lt<���s��&bj��Ԩ�����創������/����~~aQ�he�<՛D�_�/�k��-۶��=��7�����Ӵ}����$�a�������t��=kTuA	?��9h�l@M���-�($���F��LmZK߾�Qz�K��g\���LK<&X�^����c��خ�*��3�|,d�+��={��E�3< ��g�k�z/Ѝt��}45��w�=y����
*������
�}��`�Dz�P���Y�JG���`9�}U���c:�H�anh Ca�Ŋ���O����iĐ15m�A�X|�-N���Z��P�1v�uMjJ�J�)���Pk����[�?M^\�e:�lG_����`�:�ڡ�gp~x�6On[��M�P�B�!R�u�����_�l��=B{�>{����p�����T�����ȡK�=^���hÚMz�]��hǯk(SS�YW*e��Whr|L�?0�앏������d���맧���`���=*�g�E�Ξ�y�1|�Ff����궤�,��j�MαԱf�*��$�Yڈ�0�;4H�^��@�i��PQ��'�ڑ�Fڤ�҂���\��|Q�3�a�T��KD4�h�������j!y���(�4�n�R�=���S�ZR��7;������U&�~A,H�9 �����:���H䰽bJ`�.�S�T�宪	�����A�/=H�t�R�h݀�{�O[���P�hdĜ���?��q�~r?=v� ���O�l.G�:�� :�������I�W�'�h��$���Z<ϡ��pF/7�+(iT���e�:���a1�Fa��5��s�!E%�P�����4�S��C�ֲ@hpx盞nrHY��[�T(�iq�7�)Z�~��<v�S�i�:�W���2�jm�v^|�ɹ�7�m=�أ�<?p�v]�����"���sӋ�쬡|
�±�{����Evɬ�5ڞv�a���R�KtC�P�`=/��)n����:t1�H��^
���U��(���*����(4��$ma���| EOm�w��������Ǜ��I�;��ƞv� G$*�����}c )�D���]��C�S��i�B����\��A��B�N����>W������"mܸ��;F�"�u���˃l�*�~��K�N��/y��IZ��h�\�����D}�c`�0��\_�nL�7ȥ�
|q>��<|�X�5P%��y�J)��x���.�㞁��CN����kĜ��J�J���D�~Ǝ#
Ż���>�9���hM�1���)3�R1������4_�S�1ࡥ!�HöP�c��dN(�H�@D)D�d����b�5_U�����+�0]��}�"����-)��^Q���ťs�a��l�s�$��¡Mi�S&�\��"����|�6���ȃ{�ӭ/�ef-{��e��t��P3Z2�O��u��~2�H����e)](�'~�.޾�2��[��h�έ45�o�Ŝz��N��W��n^
ü	�b���H�w��6ߏ"g�-�Ԇ��XT�,�1�ׅ��1�~�<t�֭��S��:U�f �`����mV�>*�����6��ܬ��-�#��'ыn�E��Q��a�ܕ�/��a���~t��t��<o�J���<��j��(���v��eri���x�5�M�U��%����O1>�
D�'Be�y�=�E�R�m�HH~�	n�����dԓD�D����)�F �"���SF,I?/x���}v��*&�c��l�!1�V��ώS(�@ś@7��Ց�z�i#4o6��(��Ě��4�8k<CpY���y��	ڲI���<Z�� d��H�ı	$y��KS�5XP�O z�`� 1j+#��쐤dn-V����A��a�Q�k���l�6�Á��\&'�=��	����dr���,� �	�AQ֦��J"O������kM~-��sAf[����+�M��.o����@�L�����1ijj`����#bҡ+��7�#�(�"
ē 8jF�p`�:͜h�:"��+����#�C��2GS"ی�+^�3���R'PO�MZTYH)T�%�MgB�d�C
��Wm�����ϥ�6Һ)6 l��E��?#��!��-W*4S�U*
<9 M�d���¡��)���ې�!WAu�M���Q���tϽ����D�N�|�"�(�iIBߴ����5��(�2�z��*�F�V�EP��4�ɵk���`�c���d�XW��x���y�+Е�n�_<qF©+����h|b\EY�~��:&esس�Q�Y�����n���ę�nr�,���A�����*�%Z�f�⍣tn�+���j=�K�9������6Ol�ב{�:sfxFU%n���UH�_���/|�)c�����1r�o>L�vpZu$I��ͱ��kH��ψb�l�.�?Id�l�X�pd�ABL8���.�F�RZ�Q����)a(�ll�Y-�H�ܳ�F	��S�*I+}#�&E�^S~^��6o�M�MG��v�l6V���A0�h*M��a6����iBڇ@�S�&a��������b�D�V��������a� �N ΑҴ��/�<�0L���P�1L��q��L�C�(v<�&�#�Ф���O�d:��T����q)���HQ8}!Ց��&�P��T�b-a��-\��1z�0����6o-�n���2�#4՚�69s�-)-�:�9dͩc����Y��r�5�Bc ư3M�#c�4n�m]�'�? ���2��+�+) �Gtzf����y"���A|��M�;%$±��S���Ͳ����!Y{~�J�����gz~^p��>{�<YK�8z�&�F�ڎ(�;�i�X��u�'�w�*��{���?)���Mt����fw3ƹEϐ�����������Z�cN*0����#(}:v�J�C96�#��6�3B�v�ϫ��ϭб3���~K �� Mt�hf~N�6p��%����$}�K����i۶m�hӴ��y��M�ȁ��ɧ�'��P:��a��t� TJYi�@q�w��mҍVKs��W�z��04���D6+J$ `��4�l��,q�ʫ�_wdA(�'��[$ݪ\��MX�iAwM:	\���G�p��l�?�3�殍a��9l9=ۍ�1�phR(�^�U���+န	�l����4�������yr���e6P)�e8�����"'S-��7yMY�W�2H�z���&��6M�WG��� z:F�P�P2,��Q�*���%��v:� N�!OK��/9�R�$��M���?�S�\I��:J'*�'�0��g�9�t�Qq���X�]cȐQ����I�_݇\�6� K����i�rNq®䡥Q���/K��CZ�I���@�t�OI������L�Pl�]�A�CG��L4�G)�w��]��Q2wv�*6����h���!�G:�u�G8�O�»J1Ex<z��鉇��v�O<9�e�sHZ�ǆ\j�@�:=1�8��M�?y��g�i�P���� �rl�u4�ÂT�G�<D�^r��{�8�8׉CJ�о�t"�M�UjyE�-���M�	��<W�D� j6�xE҄H�#w�F�`>����iS��0G9����:��6��-ўT�W����tt�NK_����L8Cc#c<�=>G�ߟa�x��m��.c���p�zvvVt�2E��{�N�����/M2ɲi!��/�h�� �_�j���."��Ri�{iMe�=�t�*bKW`��\��a��C�p`��bO'��x�X��F�-)	�]�h\��wĹTkX��e����ث�ǉDv5�n�˴駝��i7eߣȫ�G�(c�$�$�-r\�6�'����b�A�&���j�c���x5�gl��U����vW��(<���p]�3��(f�.ge�@
���� ��4^� f�i��F�F:Ī7���NԆTa@�V�#��\G`�{����7ц�M���}��O"�%�J�c�W!��e[�X=��Q. ��%K��:6�7�N�4d	 ��٩#)>��m��:W	��f�)`;��FZ�~��~��[�����Fn����Z�h��M�������@qS�*�A�@ڱ��s���?H����drR��MA�5�&����<���*A����34�o���
mؤ�K�<@g���ܙ���b\�x�/�n����pR!��<�g���2P�F���n�S�;���O��� !�|Җa�t��x��z�����n8!H�h[��[���H�07Z �C�Rǡ\�!䨡]�s�3��dh�\�,`���Emi�*RB]ñ�n��XȈP�JEm����a�YX���y���#FsN��٤�.S�\����0{�Y��$/X�@İ���1)�w����l�.��`���<\'�*\5���B�l���5P��$�I�,FƼ����VN��7R�.,�ή�� ���i��@s��'�����P�ɛ�Lq��C!���z�F��62�����<7M,Ԟ:(���<�G1�-��@a=��i���s��=j��|~u���Q�k������ϼf�dL0��"���`��؀A20��P���jO�g�ML:�FB��:V�k7j�;�qQ:~���|!��lz�#��т54�H�b�?
�MDc�%ګr ��%;�uNI!ۦq����l�������Z�Ȃ�r�#�ը�i�D`(j6� �7H0���&:@Y��zx���z�8�c~�$GYk��4���o�M6��8��lZ[�%�2x����rO����g9l/R���|�r��i�5k'�hJ#�����9-�ii�Cgg椊���Ʃu��
���Py@5���A�(���ON�O�LP'���P
�YJ��	���p���h��N�ȗ�&2|�����<1�.��T�������G�����c�պiAѱ�)N]�m@�����W>����� 1 |Z�~����:q�SU�=�h&"S^�!3�Y
���Ԣ�Ěq�D=Qv�;O��F�=1���u����A�V�؛N�>4��s����������x'�#Vpc��;�߷���ܦy1�]�f�?Ҫ$'�9�M��17��t�Ј����k�d8��E�gO��F	�5Q�����SU�I�A.y������w�f�i��(<�F�uG�^w��`t=6�aW�ԧ󎐤YX��yaP�� A(�<��-�R��l^���H)ƕ��6���0�@�it���
�ᆔ\q�s����&�EA�˷�J���NI��h��/v�@T�����h=�K���ePM��(�����PP��;�50�H�ԋ�H6�'.c��������F���S!b���x�X^9I��ֳ�iބW�P����2G��]�65����f��^����lC��D�эR#i�ٙ��|gJUsu��U4��g�<��2�./�q:F�t�v���~���[/����&׭�\�͞jO`gG����vl��-�iblL:��d�]�-���[9�Hǎ�e�ƞ��mݺ�~t�^�,�p��$<90��[�1W	�1�9�ˀbַRdZ�|j�60[EO!s�Γ�p�qH)�����M�hrl�=��Kej�](�rmY�[����_;��B�7�|�7�<�8eY�ȳ���3pC45y�!�����hu|6��q���"������*�.�^�^�#�	��c�RG��A�&x���l$�f�P�LRp����h`�!��mś�kR$��dB���O="k��W�Y3���\�T���d���X�1V�gTeR�65`�
�;
TV�7��'�b�g?�8_�hzs�^S�P���i/�tM+&�g
�A�:S�8��n��f�*Le$1��nW;\E���LDi)���Hx��o�\+����p4���7r�R"+FFMG�`fԫw�p��
M-%��/L�\x�Xz��������B�"m�!G.6A�z6�}���A����8:���.��h�Z��1�vW��5��H_Q/�-�d�o@�o�}~�d����xVDV�Q���!�j5g9"[f��A����O?A�5�Z�s��b.���y��9���N�7����u$�]��ua�w9��.f�TH���,}�;�[_=��	�Ⱥr�
�k��6�=;MCc���
�bm��{�6nܦ��'���"mX�NsM|8p^r���dz�& ����{29�� z$����BEa��$�ԊQE���e&6ޥ}�?C�7���=�i��$;1G���ЍϾ��8h��D��J�:	7o�Js��ҬQ�X���)��[��Fk0��sU���l��8���
]�p�q� 1\W��)P�2� Ah]�sp�,X`�Њ�w�+)��P;�m�7�l�^z�~��C��b2��ꋶ/��3 o�o�B5d�[]��BJ4�X���`'s�p�_�uI�`�|�YlIո�=ޜ�k1B�����Ps��1z����&����k�E'�(D|��| @Z�<��5`4��c<�L �L�F�\ޏ�h�Fy&Q�&а�,�0��	s! �h�A[y�+Ϫ�iH1�EGh�t�A��\.jcQ��OR$vΨ �#����Q�"��S6���H]��Dpt|�bP ���O�'�����l�(�bC������9���̘_�U�Hٮ!�"%S���t������gj��#�1�]�6���0�������
e:?wTPh���8��tkl�J�i��\f�D�F��Es�Ж��b�{�Pg�m0�����$U� j�)��)�]�xa���L�4��XM eBҞb8�^���7������غQ
2�S����k���ų4�fM��%��ȱ�45�^H���;֑�ҔF4�U:!��H�H{�`�����]B7�iFTI��@��NK?�2bH!ڰ9z̑�lb��Ie*0��C'8|�}�LMq,�wLP|]��.��oS)��'S�Yt�wm�v��6'�'�ec�']���,�v/���g/�,�Z��Ŧ�f/��kK�*��V]���wDX�����!�(��؉��grv��B�J�)(�{P�mZ�g;T,�x!F�H"�	��7��$����&IB�����
�)�>'\��d�̓Gƙ�~�����}�Υ(���*I�+ukp��
Sv��2^�7��y+�"���1֟����'�����%�����,tZ�`U �O�hg�`{����E�dF�inb���6�H:!T�J�*0@|8m��@XT,�:NG/`D�E1�.Yv�(�5�_i\�Ȉ;�R��G��ѝ�½�$O����"�c�� H�Sֽ�1�Bl`�v^Fx@�gL��c�qZ(��G�kƕ��d^	� ����m�3(�͙���h,���Ru儼g�;�sj����5���/P[:a=]G�g��f��&e��K�<�t�E��?SɳL��Ʉrl7�+Bv_( s���cpp�f�Do��>q���Ѡn�<,79�a'��CQ��v�e����'h�2)�k��h;��XE#H�V=�{�k[�S�������d�ߓ�X�5r����:���#P��cp~�w�z40��g���.����P���������ʕ��P]!K7�����(�xW>_�]��,�^Q)f�:�9��6찁�HN�����NW���De@��NV�#E�Ћ�%���s9��Iz��{y�Ϗ$�,���<6��މ��eF4
�j��Ɔ��)I/M�>�I�Қ� FW��lFR�0��cr���O�.����޼Z��&����j�.�!�l���9k ��ϸ�����*JJ��tM��\���Q�Ks#�m����ET/x��J���T0<?�~'�~��A�4���з��|�����Q�a�T���qEZH=�������7�hќJ6ά�m.�<3���[2�u8g���̾6�	��2y�R�,���C���~��B����9瘒�����L��*��4d�z���k�Ɔx���jbW��*����r�$>|T������`i�f�����!]�k=������������u�W����zb��hj�e4:���D��"���d�9����̗mN��n��;X���Ҵ�.c���l6��������b�/��y��y�yt�ZM�o��F�Gg�:r���({)s�p�?go�؂��&(��p�@*^o	�J`BC��� =�c��2 *R��S�
}����@�A�I�
�m�~�x�ZY�M���<�FzI�!ՕY�&'ŋ+��Q'œ�/�|�E�C��v%�D3WWA�Nפy<�D)߲]� �b�zve����,�bl:��t+���-aS����;%�	�����B�3�jO�>E!(�O��HӋ�;�[�����X*���"Ḿ�c[�-/�����ٕm�I6�Ș��k�Q��NlP�0\՞��:�J&wK�F�4L�%VJ��m�@ˁ,�u�(ù �M\��޾�	ot�m�%�Ġ\��MA�^P�ch��O|�MBǴo�{�9��{J��]C��`myd/��kR![�u9L�gfhna�����uϺJ^��](���y!��i"Ѵc��،��?Z��F:Y �0G�%j���Of�vۊS�¦p߄��B�����������yZt�%�۞k��8�g8�ęn��Ďc�h=-`�]P|L�ɓ{١�B��`�>��wӽ��Te���l�*]y9�ʋ_H���҇����<D_����m�S�Ԩ��?gi`t3�?sPdǧvS�Y���R���"��S�A��ʦJ�ۚM�h還�z�Y�<s~��Y1��Ǟ8�޴^`>���F���2�A��{�P�9M�e6��a�A��[=�LV?��L#� ��4<�VK'��Ͳ�ch�GZ�1Ԅ����U���<h�a�:�w�Ǆ��Tຶ�3@nv�Ҹ���4��v���27:��^��#�Y�� -.֢I�g�|�=��~YT�ړ9��MQ+�@�`� lM�,D��~����?4LQ!���sv���2	��P2Ҍ��P�|B0��=�����p?xQ��H{Xca`│��d�Cғh>a\�i��9i���)gj!��?��J+l���)�Z`��Ul<���*l���Gخh��I��7F�
7J)���6���M���CUIT�{	�j��D?�b�8f<b�*E}Y:T����0Y3/���8J;���d�L���5�t������M��38J���k�(���-�]�`3�4BN'Y1m��Ro;�+��8���PX�Jh�����"agK��.`7�v�NN̖��-6�V�8�^�٪iR��>g`v�󣴖o���>��ߒ1/��쓔K���~��-��7���u��y�*XM*q��"���O��0������#'��G����s�v����|�B#cST��fU��?@�N�R�&w�-C�%�,%E���3�f��P,���=�*g�av��"�&��g�W�}�hU`���>��a5`�NLK�j.�M��'EP��
G<  ���P���Ͷ�2��K<	�ڶo�l��<l�v+��]X���_�:�9�
���>��-���`aP&Q6S�.HP7���Eі#����B��5V�R���(�xF9iIm���-cؐ�:����Bso $1�B�ʐ�b�D�*֫c���!�#����g�뛨��8#$��}���mg�/*9a��ռ]l����+"i����s}i�C��X}�n�aI�V����v5'6ږThU������PŰ��T��c- Tc�D��F��Ȱ��&j��eKn��0n���^2-�ąJ���C��m37�ƨ8��c�@��M�^ᗂ���S�oy��%�����;������1�Iu�1�^�8C�Z�F�i`p��؛Q��@�����7T����lB(R���@�V�=}�6=�D�¦1dXM�a��7RgqFY>M6%�^��?�Qc��Pm��al�ԙ%�
�"�sc��1�*k/ARN� D�SJ&֓�4�Ex����[�u�$�c�~�=o�u�&ة�RuIծƆ4�#Eܾi�Ґ�W_|���;v�������E7?��t�/���������^O��%:��T��P:�P�|�o�S'a�ҫ�o854�Uf�yQ.x~q�*��(�u���r�ku:��,��F�M'�H!9J����� �6�Y��:앃�,�S"��꒴�'BOw´𫰁Ǧ�U]��F4 �	���װ�SO�˃��Qd� �KX�H�O9dL+0����DS<�gϝ̉�BC�>ق#���F(�L�����A�=��<�8##CMT�i���zj��'�i)��|e��4jy�:�!�Td�Ȼ�.ĞS�ڂ+d6�=�S����5�CZ���9�	)J�6m��D�D*�)��E��]
>&Ol˺֟�Y(�/*�i٨�V{�r>�h��t�^��$�U`��7j��I[V�0�NO�!q�M<(�_ʍ�g��V�$	c�M)X�A���x�x��	M�G,Z���C�|I�a���a:&-��6� r*j6~/J��C�dLQN8$өg��4c�+w�Z�*�c�v���S>[����/�I�gs�>�8'�@td��A�N��
�����vPJ����¦o#���)"M��e�BE�D�e�����PM>9��"N��pM�h����rV��S,��)�X�Z�n���<�LSwD|79�/jW�ł4�hG(�@�X���-��3�uz�;ibr�*e�z9�4P0������D�B�=�2����ڼq��/�O}������>*�2���A���פ�b��6�z���td��\^&���d(��[���B���о'��ĚI݉yrU��6><2.��\��ye6[YQ�I}�L�Bn�Z�e��H{*��<��I�9���!a<C.�0&�B�A����;0��"$"~��@@����EAԌc�Z���a^��laH`H�3����ʲp<W�:R�:��2���G���"�Bz����4�"e�K�ׇ�r(T,/����
�e�:�XmyN�VC^`^��τ'Qݓ&��
�Fr۔�˼������j��
�sb��'UW+��+� @�}L�/� �z�V�[�<�n�6��]dIĉ�#�-�bS�JsC��oSQ�A|H;�8b�^��a��N��_�dAO� {�{��5j}���[�r��_���r��&w.�о�sh_�)>���#C�>��%,� ����g`68c��κ��ӱ��M�!��+������K��#�!�����y�0]$���o�J�ϟ�4?�@[�l� Qx���M��h!ұ����%���V��;����^��A��7��T%RT���fJd�2�2ɨC=m��˴#IW@Q���_ũ��'er��;D�u�w���-�i��x@��
C����e��s%��V$*��E7�ࠦcҩJW����r� zrŀ�B�hK*T.���uk�ѻ�����8:��1��}��_v=-4��޲�@������o����5�[p�@�Aa�=�R���-�/�!�����۴}�zz��?@K<!�o^K��hA�3�'��EJ��t��I4��;���n��}�vz������o�����H���;Eŉ
=s�Et�O�_}�����w�v����=T7�+5����ћ�ܮ+�'�y��𕶍HB���{aG��9ɞoF��]8KW\����a��L�qD䷸4G�c�H$ܭ�����?�=��[����{�
���C۸Ɇ�΋&d��ڐ-s����SmiE�=f���c�Y#'U�^�f�l�k��20%��&��U��(�^�np�]�'�t�Zh�u{�ۗ�-�B�|T�KG�SH R�3�&[4LE�~&e�tJ(F<2z� ��� ��	�=��J2�����Cai	NeC�F�Z1!���^�ɚԀ��"ck����pΤd�=�p�8M�0�0)l�h�B134�:����E׀B���r��bb��ZS�AY�P5�0>ұis����ʫ��v�mw��2�t(ʻ�H�
)~��
a���Bjdx`@rە�v(W*Eu��,¾���=�϶�B������Șwh=�b�V�@�|KR���H���99'NE%��M��T�A6�8-��Y�� \��^� ,RĦ`(n��� E�pV����.9X��񥗬�믻EB�r�ɳ\��3�yK6<W@�!�}%�׍�o�-�n�8&�Ʃ�d/�<H�ֲ��9����ԆIJ����T.>�fx�}��CW_��}|}��{8Twi`d���U�]浯z��׮���t@�F��<|� ��=亂n��zC����{� ���S�������|��t�7�/�vڶe�~|/�f��?~����Џ�� }�ߍD��REs���B���6��.b���QBY{:�ҸF�o��.)�%�3GS��P�^�ڗ�g>�5Z�n��Ο氱�u<�}ZZX���������k���sgUr�d�vl_C���/���7Q�!:ql����jBdtأ���Vzލ�������O?M�����_���}��Y���T����]��o~��ż������ۑo�g�!�坙=d�YJQ�L�)�RI^_��|a%�|�T�]C��*���4�D�߶���ה��jǙ��(Ǝ�]/Z?��\%�i��lL��kXk��d:�\C�吥t��X&gM�#��]S�����3��Q�`��d��\�ӥk����'�'�}^E�CD��^��(�����I�� G��d@��qj�F�;k?���ƅ��W��{G��� b洇7޴�(�����"��٬�3�w�є�'cN�ُ�et��I5���h�xQ�@�Z�1��SOE$���E�f��y��M@q���c�)0�����H�id�E))��vcAi\���o �>�[��iM0r�ّ�ntd-m��M7\#�������\�l*r*�~��v�D�Zs���g��^�cz�����ϻ��Uy|Z�)�����M��o���s�5l�������|�|�}�M�����{�,��D������,m޸��!��0ϋtR�o>�^zݛ~Oh){d�=�.mڔ���Rz�K.��ܺ�L�\�Nz�[>$8El���m7R�]׽����i��G/����eZ���Q!����M����s�LQ�ӡ���m�8d���ە"�Ml]�)_9��L�Y]K�oJ��ԟ
%�?�G
D/x�#�!ڭ*��m@������R���~�w>ϋ�N�y���������_��^����_�	{�|>���7^}����[o�F7]�W�ڗ��#��e/��zp��	�Y�h��Y<���sb���$uxN�ًo�����M�o��!�e��{�����N��0�^B�=Ú�]�g��$T/�1�90�Y�(����p�.$};j>�*O<��M#��)���;�M�.0dO����K\t��`{Hf�/׉�dr��=�`�*O:Z��\�ߏa|�<�R��W�*B+_�(�o\�T�M�ؤ�]�M�^�IOEnh!E� խAM���IC\X��B3��J6t���ܗ+|9=�8�z�Toh�'dϕF6�U�p� �j��ʈ��L�ى��C���g#� �64%�����2uǵ��$)K�Y�8ZMJ�Y�F�(�.j�w5��`��-9V^�5�a��GZP��Y�/}���%\����f!�E��|P&�iee��}�|nh0�QK=��C�NfOJF� J�u�����C1,��_K�#�N�N���T�8GB�N�׼O��G���9J���W�_�l2H3����}����X�C��w��r����F��>v;ا��zכ��ʂ���s��^�z
[9ʍT(�}�o(��Lh(�Xg{>p�n�q��\4N����ruF&��9�{�iI7t�Р(ݴ��T$�X[�����<b�t������I���9� a����n��������MDD{�<]s��(l7��w�9����"�Q2�R���7�k_���?��W����vC䱭�����i	���oߥO}��40H"��1򛯼�y��O�ϻw]A���s���t˵�����)K�f�wl�����K���� i�e��А{<D�=vprK���^`�ǸkO�;�ø�cS!������O�`g�AA�X �"O����c�k!�T>�I�6Lz6��B�pV[��	R�߄>��\�S^,z,ߐج�]���q�5�ɶw�8_��\�^�������I#�s詑4)v������ע?��u(���F��}��O�v�asC�.�5r�£m
�H۴xBu�P6�*е,褮��9(RAy�G�� �udX�6�#60���m��3��V�F�Э񕔥�FX�}��C�S������L�� x��m�W�QZrӖ.HW�IhfJ��DJ:6.��т�yQ�]ںy�7���r�_��M�� ��Ԕ�� �I:T�rx��r�
C��b�z��A#����Ō�K�����*x�R
;9C����ŷ^O�~���[������i6>k����e�m���������c�}�n�_�q���"��>Ue��?�[t����_qP���P)���lͱ����}2z����{�?���weBhWj!�X���2���ӑ��C��7�B~�F*��#�V�|�)����7]���d�kV�uxdx��Ϝ��F�zBXx�m��9��Z���`']r��x����7���5Mn�>����=�[~p��?N?�w���-�/���dEf��+O��Ǐ�_~��鵯�%z�k/����O���}����ݟ���2E����E�����<�po��׫�482&q�fH�t��l��;` �Q����.���5��0����E��e�����d�Q+ʫM:nĴ�J@ �=��,�(�&��QA��^2���,�T!+b�j(cT��5w���t�F�MQ�y�az�<E���c�%�=D���M<�zbpƩ�t�J!�1✎Ұ
]��J[�nhx.�I���1V���"�wlRL�a�4ߜ���F��Q����vS�F�ɥ�	�z�����)�d���2���[u����?"$^�(����
�~�s�t�:%���9��B)��íi3��&r��e�O�٘E�[o�����f/�)@����E@���v���˥�GƗӏ~�0��R4&�\JI��+�*
o��=+�N�n��c��7��2l=C���m����h���Ŷ�A��G��w��R9KgO��o~U����?�����ր���^�����7�OAz�reZZj�%;7��9x�n��9�O_��[���y��G�D?��b�g3��m(j�[��#�%u���d�$���/�o}�5����2_=A+Kzɋ�JϾz�Ο��}��t�5[i��&�V��.���k_��,*�&bz��S���x97?#���g������ �}��u�vt���yz|a����b�-W�U�x�]GQ^l'�;�	ڻ��v~�Jk�JJ�k&���H��p=p�A��_!͜���z<�:�y�\����k.�m�r���n��窴i� �� 1����O�=��	y� �ٹ3C��Sex=u��i*����T��Fw/�tl"�� �.�>�@w��`��?�H$����@�FD;Z�[�/�b�b9�)QFQ�M� ��{I�:�]h�fqܧ�8�n��t�&7�)çy��g�IKm�*���N�U�`c,S�S��vD��t*ڤ�3}`��;�oDF&Wm��}:kZ����X,�}��ύ��_)�����t�1�N[�=IMh�����	C�P6�]o�.DZ�_�3�{�ь��u�D�ٌs�z��J='��H!����b����g�f��&=��g9A�j��2ŉᐡ�&�SIaD?�C���w�y�Eo��3�rF̻T�H�f��+E!�+�T�ѣ��+��J����y΍�鹩h��f�ݡ h�Y'�@q@�؜}��}������d�=1=C�<�������(-��$Q~����n����'��(]����3/�����:��g�K���	�F���zӛo%��v�XO�?���5��^���_���s_�(�4??K�kI5-��ߥ7��U򙜣!�>s���JT(�ϟ�0������ϒ���7/���J�س���"�pW��هi˖�0����tB�.�P:�'�Y)�e������ٳ�����Y�6Ŭ�i����m����o���i�z<]���< �b�n��b���M�go�����_F_��]�m-ӻ~�VZmO8(�Pq���:t�]u��G�K��� ������w��hqѡ|�8�'F���s���Q��G������p��tӥ��h�7�x�fk.?�qYx`nS�SJ�*ȧiq�Q��0����lHn<�0.�ɢ��.�5X\e�Є��#4Z���pq�6c��ܱ�U�f9$Vs���L�xH�)7K`r�6nSI�>���yl�ȉBh۬�t�u��n�w��p2_�p��'A��k��zo�.���l�̽��B)���� O<�C+ke�$0��Ѿ�r���H��6���3�>0��T,䵵�TMG����yke4ㄈ$�F4m.�>��J,4��+�t��-4	�X,\(y��
,�GL�ۂ9-K�7��E�3�Pd���������(��M��qQDO�m������G�p�+��@�P��_3F�6NҦ�i�����Y�l��JrFɏ6��;���f Ă�VGy=�=�19Iw=8Ǜ�6�>����^�\z�KJb$^��п������
�}�_��^��װ���oz1]q�U���|�on��}ڶf��}��O�����b@������?��������w��҅�<�����/���ˏI�L��o�ƫ��d4@�k�$�?x�n~�f�������ڱ�H�����/�O�N?��!��YC���g�o�* Nh��uX��Ɓ|9��e��ٰ�7J�s�����������7o������)���6KN�[���=}Z6�t�v��D�汔�¯?y�J_��7���M������|��d=�����	���ڸ~��>z�/��=�Q��:zb�&��h�%���ctˋ�K�\���M�O���|�f�K7<�=�g'5j���g�'��#���*O��@��(}5�c�ϭ�0��f�Y���N�Q�p>�c[Ń�8:5b�cCv�jǞ��h����6�nU���<4�EkDl�+��3ND&$9l��|u�zZ�����yg��f�M1�jH`��S67�
� �OxQ�m9�&�F;1�flzX���UhZ�����D�}�������H~��j%�g2��#�e��4�i���Sg���")ƚ�	����H�Y����r���q����lm���=9Yճ�l�U\�H����n�Q_I�����/���Q�����n����ܱ�52wL�5ed�B���m~�pYX�qa�iL��y7:�lx#ʛ���ZH��ĉ�=ں�5t��(�$,uD37^�&�B�0Qb>���=�y��Px�t˥;�{{���Z�R��u���?�﯐�ڰ!G�7��_�g�����J�n����7�9���,�#�Ӄw�4�y�K����<k7=�Г��?x��O�m��D���;�W^�rZ3�V��%6���G������A�`M�񆿢�'���D����7�Iw���>�y�>���T�T�h-����n��?}�n����/�A?{���2�JA&�e#۔�T��@k*�j,7D\��\�F-��|�_ӗ��NtX�x��������x��_{��ө��[_nYY]��x�Ûk�B�BD0������ح�D��:���4��gMbMD��qjM@Em%&�EFQ@����GUQU�����g�^k��އ����xu߽�������Z�xP�$��o�I��hJ��/��r�^�??$��5�}�I���{�P_���'�����/��ծ\|Ʌ�zMȓGNȮ�6˩�����y9�����c��e�~?��6�@[�����^z�,/���8O��]ߧ?�zy�5��{��C�"u���Er���v�
�i�a�#nby��W�^K����'|H��:�����8 �ᘇۛ�s�ǓGρ�A��[bGJ\�/�z�!(������A1\E��<+t��y@�K6$��ů���w	�C]3#�sf��)
����ׇ�)`��=9d�3ξ���b{�O��q�ڐ�'�ŉY���o!d�sV��th�P��}B:|�l<e�t�m��y������ʲAbi��<���3}������3�UL ��3�u?r���!����G��E��0a��[i��Q��˲<���Xd]���� 0-�W �#�eP,�4���@��wV��68�����}s"�g��bW^���h���i�znJ]���fؼ�t5>8�!C�ᚤ� 
���֚|�Qk/hpv��O����\����'���s�/{���qK��z�U�����ز��$!O�BW��J���c{Vg�~�\��/KU��������u�E�����ڸ�9�T���ꫯ�#� ���o��89z__����B�-܋�T� ���2���_�"9����/x��\�䁟�э�Q\k�T���u~qC���kh��Xc���Ǳ|�{�5���u�"[���ۗ���=�"+�/��by��X�A��/�+O�Yg�.��E���>�v���~K�;*o~��K_��>�D������r��~ڴ<1ےgԥR�-{��=�匊�u�M~����q��=�������21S��2����{��}c�N�f�0��̔���ϑW�΅r���c-\��Ñ��)#k�bl��I:���u��+ʨ�"S"����2�r)y	���^�ꦭ�I��fy�Lf��.C8g�1?��UĄ�A��N>m}�Sm�#+�Ds�#&$�9��P�p��*��K�{����h�tȦ��+I@m;s�$t��6EX�b��\8��W!�G��p�:B�~n���- Uq9�D����%���09��������m����OU���%f�q��J#����S:c�Q��d��SJ��Ͷ��0�]��X����k�7�m`�k����86���������|�a�ϼ�������Q��q�to�_��[�+�-K���Ĵ�
�����wك:�j���"sg�m�W
�G��uHg1���5�-1��`�}�3ܞ���_Do�)�7ѐף��De���y������>9���wMn�cz�\��I���xp�z�k�ؑc�xw�:MN��4�`�Q��k���s�&y��9��gn���E�?w������r���B����ʙ�\�)�^��~̋���?�m�#����o�U/��<>{H����S��]����u�l�f@��9_E��/�~�|�o}����|G7�@7rM���TH�:���x�Q(�����b�^����S偟<�n����"ټQ�1>!�fC���z�F17���ؾY��o�5��eӖX�w����w�L��pU��Wn���A�w���}�f>��L����WK{�%S[D(�u˔:��n���k&����r�����'��#����Y����Ck2Q��u����Y;����J4iT_���CW�px�u�:6�F^��j<9�Qr�$�>��r�eXY�q��*��<��R"Lm0��#rB�.��"��G��6\S֜9��=��<�#~o�IE�]��B���E 0�� 2�w6`p�+S6+����(��� R��}~�S�n�.4'��@��yC��e��V�K�.wlB̊`=s�]G��5�P�pd��,�{�������I���C?�瞱{����O#��_}��F����7�GB�6XN+A�:Gҳ؞���ށyc�(s��+�~@��񄰤A��:�:4 #��"0�^������{>�p�=6�Ǫ!'s2i���MV�!ǉ�(������?J�K-}|tU�:�t:��Ѩ��yUh�T�ʌ��s�%ʢ��h�z����c׮�IK�S3$��厽��������{cf�1���7ɑϕ�c�F�-���M���E�7�X�{���cc[%V��a\������?'����ո�聇eaa^��� ���w����
��3ٰ%�O~����]+W��]�������BwI&��L��|X�fx����\�iߜ�ڊnwO���ڹCf�jr�����k4����z�:DZ�WJ��%+4�R����l��������w�_�׾���O~�52����1��ujJ���~�<��|Nv�U�����R�d��@��_��o;(�>7��wR>��o�7��{5�׵�@Hc�"��#��}���~�<��B�N6o��go*Q^pٳeu���}w��֒x4h�rσ�2���ɮ�Dc�	�e4Y����]����dM�ˈ�Qt�.:��+k��d�d���0����S��?+�Ad�� ���8nNq-�@�BPֺM�H��"�Ͽ�!!R��_)`�p��x3fn��V�K�)�]t_�Z8T�R�5ψ��_����1h�Ǵ!K��ֲ���Z/d�Y�hBZZ^/���I�a�aTh�Ր��>��pʶO'A���	 �6!��\[���g���@<>��$��M����%��?���܃�x����EC%���k�ְ��[/0l����$�r~n�6Ni���lg =�	:�D�7`���lE3�n�?Ugd2ħ�5�\��yVJ�A.=W=S����d��P�W����zvϹ��q���=��D�����_y�VF�k]O4���0]�b���w(�^ėr.�&AM�.�ٞ���ڮA��;�冽��M�xQ>������/~�<yr �����U������\��u�I	�U#Hw��9y�U/�Rz{�����;�ɘ���_�5ӭ���¡�x���9g�G��g���$��m��g���o�׿�]�z�T���,�}�K?�W��&]r9��3����gr�wHeԇ�F���.�1��w�I��H]'�(}��Gj�?}�M�}V����Q������"ޣF����u������|���HuLdv��l���M���a��J��AA��g�ȥϾZ�KC�,ʓ���7�{>x�'���,f�|��_�,�er�K.��,���h8�˳�?Gn��~M�')�koN�I�ړ����i��Z����2e㬴�=���������|wXro��u�`������!F���u�=���H��b��΍@("n�j���b�E��u���G�J��j��g@0<U=�,�Ȱ��Af��q.�u@>sW�����2��uj7�7t`��戡�96@�Y��Yᵞ��Ű�<�~�v��(���?7}�Ԅ�[x52�8 �8d���a�a����C�S��9C�Fk���Q��<٨�f�.y�s�L�x��;'Q��\?�zM#�a<l8�e�y��^8�
B�20�Y���w����|+Qbn�(I͈�YR�3p{�ܣeܬw�GחīJ��s�Q*�'�	|�e�"�)Z'��́�;�ەӱ�����M</�&�� �.ҳ��O�.ˁ�;��O�K.������.4�{{�i���|��=W�εX�%'���Uج�ا+��9{�Y(�^�ZQ��v( �pu~S>��/��.��/|�5/�e0��ab���rr�y��<9D�~�[ߓ߹�R�������k�ڤ���R[|��'`��MSݢ)E]�@0d��	�Ls<�o>~�|军�C	�bA�x�.r"��o�h/"8>r���_yX~�W/��=�j�Kj���Q��|�T�D��р��h֤�:&ͱi��+�,���u��^yn�6~�����k_~P���o��]���-�|��;�����&��E׊_�H���?����g�Ot���o�[��'o��\2-Om��_������q�&o}���z��+c���iˎ��e![��@3���i	I'�఑�B|8��[-���6��dlb1e��Y����A�H��F�[*9�(e}���'WFx���>�U�QV���A"?�ͣ�a}:�o]C�D��Ĩ)�;���u�y=��$Iī	�������'�E�,-���+p��,��>˱h���|c���l]�ΡeJ^�ƱK���4�PE�"�R	���K�%w���y��9z�<2�Ya�8�$ #�Ʌ��d ���>��g1B�h��3�u�Q
/�H��~=Ϝ|�Np�A<Y���W�NE��1�14�a���T��\�;"E��)X8
4�����\�������	x6�a�$���}�Ig}8aj@���>��G=B�8r�Q�1L=r^��8>#��9����N�k��	|G=_�͂����j��5�h����5�����j_b!���]X�BZiU�(��t}
�����a<����-�I�|�m,�y��jcr���	�������>|���U���M�4�"��s��އ�#�����@�?�|~�C��%y��&�N;U��Rj�I����C�/�3�L�A<�����1.a�E�y���o>�JF��K"w�s����o|P^������YT�����e�y�ȡ����������y��k��2����ݥ68�����Ҍk;l 45�<�ȥgQQ`$�5=Uu����G5��,����2^��+E�>�"��Q�&��ZR�x��&z�����ٴcL4I�ݧ�"?���}Cv����_pnC�#�����ƛ����ߔ/z{ؿ�)en�����)���%[;*�7���#��fY��K/^�p:�dP�A˄ȷ����S|8�.�Hs3t��{�p�j�(.���H*�$�JYΰ�\?@`Č�&�f������0#N���������"�� !!ב�_덷�ԣ)e]���J4�m���`����̹La���P>�šD���m�CT�U�3Ǔm�S����[�����y�������u:�6^�>+4�RK��.����F��IX/&E�T����!`��B.�\;б��s=)K�$F��n���54�q%`��5�P4�Y�-LT���F^��EC�A��_P	��5|G��+�[ ̙;�#�6Q�w�w��F,�H���v�U5RDq�4c���|2����I�T�6I11�>k� !f�4���vl`=��B(���CS�p*��!�?&yEת�{C��4�����\�={�ڵX6N���b9y2��C�r�Eh�W��g5�����x۪<��ͺ�v?�y�	Y�Y��U�ve��Tᵺ�g�x����m������ ����X�<}9�7n�$kk���Ƃ�-�3�ȣ���S���\��-4�W�����i[��)7|�r��23i����RٸG=pT6o�&/�g�Mo�B��C_翿�yϐ���?J}j��/<"���d��iY>2��CU^���z����%��䊜lo�Mg]"KO�J���5� �D͕Fľ�>�e2	����i�U�����Ɂ|響���J�˿�U�n�)���Y\����,�9.��t���hj��6��������^H�쟾�Jy�U��쉖l�N����'y�{_%�|����.�T��ѣ���s��?��x����}��r���������{������QШ6����z���pW�ա~�CKc�jԾ�OӘ�����M�^ӜF:+ ͪkj��$�.RQ��4�����DIe'��c-�e����L�φ�pz}��|_�zz�!�Qy't�S9C(��Æ�}1��rL�(84�ʡ1��BZCq�&���&��}��jŹWr�GCtB�c�]ҡd�'�+	]!�0�0���δX�������!���3GY�uq��!J�0�U,�y&l9F�����v+��BtB��2��;k2wrM&&�R������F][RSG�ʘ%3��@ɊZ���GY���ؒ;���NXC�:\27�Y<SC���3�(Cu15Јh6+��A�).�j������.��{�kal܏�j!�m�xkB�����Ƨ뇞Q-���5�а���C�s�@�٨�h�m��0��0�>�cK��;	����N?uF~���~n�C�}�p&��>�!�w^��4��<��Џ-�D�)i��,uӍDֺ-�*��@[DQ�FY�ޔ��z�>y�p������/0�ծ�Ɔ��}�	��.���B���Qy�{n���y���(�^��ĸ֐��cyɋ/�n�7aT�îS�ȱ���5﹉lt�^E~��A�z���_��D"���i.�y�9��n���8���4��s�EDQ!	��Kֹ�bh=g6P�0�PM}j>�k'Wȥ}|~���W��z�s�y��'�w_�>�D������@��iv��?�O_:��|L^��G�W��uP��
��<yt �}��2����g7�=N�����k�� o��er��o�H����y�Y����t ��F�4+�b��zE��*�����T�������o�&�^�����a�5���QECNꐵ�دI9���1��V�O�\�5�q���)�������E�&��و�Y_��A��3r㾙�������|X/r��6�_�{�E��!:Jn�R �Ӡ��!�"X�w�rz4��[�9�*xp�r �{26��lk4j��1�I	�݃�ȍ ҵ�����N)�pF��~േ�,�>�����0�0�2B_��H Uʌ�H`l"�\�!�x:}��k̯��L�F_��jSz���oL�p��,s� ���X���P�}�,`��2��G�������7��E'[��0����x��)�0��S#��밍�V�����"x��ld�m>��齗0Q<�j�Р+fY��2?�bc�d��N�jՄ��p(���id״��Z]���|"g���ز��yM�29m�~��-���(��{��HzU��f�d�'d5��ܺf@]I$��XS�X�0��R������&�ov�E�m����ɉ�j������L�8�lw���7ccޏ>qL������Lt��	���7���ކ:��|��BZ����{;D�S[��%2{�d��ޘ NO������|���5��B�R�ln�迥��ь���+�j���3�6�{C�OLw��EZ��0�H��cS��4��Ȃ�}wA�:ޓ��}�z;]/��cU����Y[�QU�P�����'ߦFbN�긾�V����Hts�42f8��m����N������8��e��}�V}�/����w��u4�����k*�ׇ
�]���W�%�h�2zf����9�9�P�P�O��;j�$t�����!��pc��ͣ����f�O)E��I�q*<ؑA���V妱B�׳�eQD�D��l+Ox�F�F<��ʇj�d�1�c�jN�i�Lr�8�?��$�2\���N�<�0��`�+����t�#�o΁B'рŘP��Pa�����C��C��b|�&>���ȖA�ϫ8R�QS�����gPH	%����R����� �9�٫��H�5n��t��5�z����̺�OOMɂ��k��}Ӌ���9ҩ �<B�[8؄��%�I�rs4EP�>��~fQ\ec�8�C:k����S�,N�e�a���@0F��s]�(v��cڜ. ��8dd�U��pm�=���&{�kD�B�sq�!'L�cCSm�v����e��>��0��j`{���"ep;�k�;~��Ò�sn��-RY�}~ۃsB�n������
�PC�Hw���E	������'���9%�pLz�ey�DS6nڬ�.�wB�YJ:N�"A&�̓�3rx1�ūӈV�!��>.0�?�ex���K��v�>�K/!v@Li���!�t�>��P�̔���RCu���,,.ꦂ����a�k`�8�&alnr	�T-]PA�Z'7�6l���F��s���2=��������z t�4�N�c�PZ҈��Fk�1�$�8��E&g6�E�k�i�N���,--K�ڐ��Eٰi'�?�;j��q�Ν�e|b�)1wRvq�S���8M}x��U�j�N���Kx�h��*w�����Q�!"��\5<�g�ˍ[N�e��|7�G�qH�W��[Iu�u'N�XF�ȀX��y��Q5<��t]{?c}��w���φUK;D^04ތ�r3�C)1���B��چ(-�p� D��4R����9G �L|?��m�e�'�����l�ˎ���9�0Թi��آ^5.�$#j8�棁��)�@������{���9��=O�s�p烾}�Y(�	x�%>�������S��=v��[ZK+�87��$Qj�Gt��ğ�I͠��]70"����g���4���q��5���[,0��}�&p:��Ǽ{5�痋�п'�%B��0�F�F6R��o�W5P�ꚪJ2 �GX��ñV��L�V��D�Q�2��`f��'S�� Ǧz��[��YV�V��{	��,t�xj0q� �_�K3c��������r�˪+��M[���|�g�,E�X����6�d\7FKmh�K��DK=nkD��"�R��.��B��,]�K��R�h��m�B���f%CF�՘ng��w�6�.��{65U�p3V#+�S������4��wѽ���46��R*.�)" �c�G�}�d�tk������Gg��j��5�h�<B���^�M�v��͢j2��6\XQ^K���L#��j4F(�T6�H#r�,E��Z���T�}�g����j�a4��]Ҩ�d�:�Q��[_u������yU*y�� Y�	S���X�V���W��&�YW�s��x�HWs�萖���t8$��4��P+*�g�Q�����fM5�@ X���K`�Beb7�^y`�-4�P���ZḨ���hH�����a>[��zՔ���C�����+v��"�8&��^���5��:�DŸ��]��@�U"����%��j|����rW��x8���!%)��ˀX���������-8E��h���DA�˱n�,q���MX��:N)��u^D���^�0ѵ� h�4d�͚s��@H���]#[Cp��j��&�S�v!��o�tɇǰ��&��ք|�s�0���>�v<C��'�з�c�vF���u�{�>Tx������S����ا�#]�>�y���='d\~íF��OǙF��V�y"��  -L�1(��!��'�V����S^��p�+M5�	JSjOj�Zb�E�Ȑ@VQ�4�٬MjuڬH�{g��|�wL�@]��]{&l  �IDAT�C��MnN0Pu�6.�i5w��ye��&7��U�4#DM�׸��x��لEs*�� �u��#�z��	��U�T��@���;mM+�����7t��5���Y�\`� T05%D�O��3��4MF+r����,�$��j˶�u������2@sb~�6���Z��k���8��v�憪C/l3j�Yk*gb!�'wQ'��n���ܸ�����ߨ!WB2�u}��)	,i��z�0�C�ZA�(��g��3�a�\�=eY	�>��� -�\
(s��@^e�?^`����bpDP���s���8HL�b�p�/-�:�ȱ�eY�I����P_ѐ=:/0��@�!���H�<7i)sT�S���(ע��Wa�m�!�G��p�"!�~���I0>>!�t؈u�g;:��a�+�ny� �-��}
�A's��ꍤ.ݬ�g�A��K�<��@��:"��E#d(>���#��}�7�Zf�&v�eD}F��8��5�gT�O�3Љ�C8�(�z֌��6�c�"�+�Dq�l�#u�-�B|D����*��� H��6֎:�2ԺR|�/J��-Q�+�jӚ٭,򘅇p�b�'�>�1��ȭ�3�hGh�i�J/��+�+	q8�D}�gV�x��B���}�ɹ6�]+R��;ę�c���r6J7�f	�3I���A��K�aoE7*����W�Q���g��F��ܠ��#4�����#��DJ#iM��h��0�p�A�J ;w��!IH�S�&��*e�Z���m��؊��lL]���.�7��.��ő�d�cc>��74j5W��-�.ܨ)�"U5(�1Έ�*�Ho6�UV)@�F~����FTO��4(����5όͭ�w�u6�.�A��i��&�Q7j5�(o���8SC��s|�N� ]4a�O8��F�Y�i��(p��O��2��s�}�at����S�&�]1�`��a��&��&�B�k�$\��&vI��&��tSq(�U��L�u�"�"��H\jV����S4�=1��d�p��~�z e$!�Az�N�(�\��<|�:-S��=�sRLy��9Ş�>Hp�&� FY÷I@��Ф=w�MF��k��Q#�G�$/����g+Q��IF�F:�F�`�o%/:!7��ʎf0c�&S|�Qg�c�L�.r�ʡ��2/B�� �MG������:������ڱf���Z�_߁ֱߣН�"�f��l�ו!:k�B���Xq ��NfnMLl+��{4�ߴ�g�A�2�&T�d��4�%3�X8�*�_���[։`4����IX�w���;��3�<UZ��2�E���5�&W�� ����WVИ��똄�3�����"�4x��� [�Y�&	z��4���w!���W��R �*d�4��^u�a��R!?���(��}Dό���O�,N؀><�,´iD3rUF��\<��:��M��dZ�)=p>&��]]�ծ����s������
h�iJbS�ʆ�R������0*H�PCw�xm���A��-x�&QA�.Y��~�#�S�0�ZkL�2�t�!b���馨iQe:���vrw=|�8�m���,'�j�����N��q]{�0�t�ٌ�9a��mk`���ƌGiJ)/�����n�����C.�.��4�"���?��O���D��	F�t��h�&Q����[#'�H���d�~H���8<0��R���j�%,66d�Jy_�0�y1Ԃ�`P@���1hP`}�ȩ¤�7�����NaA�p�0�J�0�٘'e=ɐ)�J����1#O�ؔ�aC�m�	�1�@J��Qq�=d�`���2D�)��"MH�u;k�K2�7i=�o�o@�8�����b�_�s����2upOC\���9��Jٲ���l������ܓY�$���1xD�l��S���q��%�y_��Zl�P�([��<��|z	ݤ/}���1��ם�#�a��)�����Zj�@�V��������j���C8bD�N��Y��͵��KW��i���׿@���z/��8w�b�fe@V+�F K�]j�]u�������iu�c}Hm_���1�B�f
YZU����Dg=�hLԚ��J���J1�&���j`0�Hw�Ui
et�z1~�jS0��:YM���НUw��P���k�.�k�K,#����Q�PX�+����%���ҳ4Jj��� n6O�4�J@vKTT�L�T���x��L#��?b�Á��F5��}o��6D�t��lH *���XUS{X�dL#���8]:��,Vu }���+�Aj��)3�~ǣho��Hpe��	9������"�aeE����7u ��s(� �z�<�L���B��jXFP��9���p��0�d�C0�,?�Pbu�H�YL�_Mf������3��c�H��[���.JG	������y�W5���t���o]�W�kh\F�^C�FpS�e���������R�%!�}��&֋1�o�鞀�|��Ҋu.��mY�_^��)�Y8(i����^��o�x���K!ZF��i��Ȍ*4f)����w�>p��k�o�D��|Ei�R���|�pV�5rSD	?~�s���j�֙(���2�'�Bݶ�i��i���+��>HIt��zv�@� g �Y&u�踐aFxް��t&���9;D�yf耕�Ԍ4���B�y5+V�;)�!�����4�A���8�_�:�1��#�L���9��l�w0���^O7Ky�����pLƧ6s�������Uf.Q}���͢�>q��vD �e4;66���%�e�����8�D�Ζ�'nJ"k�}ʗ�v��_������"�K�bƣ    IEND�B`�PK   ���X����7  �  /   images/2b66d102-ef9e-4dde-8ee7-817842500f7b.png�XwPS��� R���PBU�!��B	M@E)R tH�J�^�JGH�.ҋ�PD�@QJ	
�}��͛�����:{�{�:���={�8c]����dddtp=��YD��
p6z�d�>��zh226�s���v�^"������dTg	�E2�3v����3 �)������7?�s��ܒ�G��/�?�مg��EAFv�o�{�/�}yU��..��=��} �����ɋ	�F��>/��-+�>�1�Z�%��|�����p%��9�#|*xPݎC��S<�'���o�9�^>�W1L�Q3����.�Q��Օ_||�*~d �֋��'uy��j.��9Z�*� �u��+�>E�� �U�L�.5!>�n���f��f�q�7Q�>��-g�_�T,�X_k����>�:�c;����F+��g?���r�q�1�����Uʰ���r�S[0'H0]l��?�הۖrm��O�������98��W�8
�}�)��;C��r��3���&��?�.���d��ƛ�d��M��X�2U:B�72���/l�b��!�#8����G��d�{��x���m������#럀�(����ū�e��}��� }�g�
�B�!��R�����R��QD��z�_/�)��1@�2���X�L�d �IQ�l���Fb� ��yg�W�o��t�Cy =�(/O2I)IGP�yYr����?"yd�{n�y�kΊI���;���!����jx{����QB�
�����8/�<$���9_�B{���H��w���;�a���S����!EK��ű���"���l�4kf�Z����Y�5h[Y���z�_Q59:�eɔ��5
�Iu��qV}��Ԕ��� ����TH��.���F���b�	�mM@&�cA��	�)�����mگ��wD��M]�_����Z�)"�P��R3���Õ�m��~�y� ���,[=lo��� ��8,�Lć5��63�*(L|�H�	�A8h-����"Ҍ*{D��e`ß�Cy ��g\.�PK���$CX���U����a0|�.Ȣo����G��EE���Ϟ1�$��|�B�ܵ[֘hkת���(k
E=��/��-,�$bb�MLc�虅�/�6R=xW��4����ZЋ'R�Uf�8n$Ⲷ���5]P�I1ِݰ�C�d��{I��M�7��B�!�P%�A�ml�A��ƀ��$�R�zi�pT$5h��h�p�V+d��<�~`pn�Ȋ����	@7=*谭��x8-	�v�'4k�߲t�]�Eo��ʍ���\~5c�U��-�Y�Ԅ ���D���҇ӌT�L�%�I<�X�(�,v����Wn��L4����P69����'8�r�rI(�d���`�G0�G�14�k�:���
��$(�;���lEo�y�B��^z. Ul����i��n?	���L�{���S�1'�:����\ϴj����^P".�� �]�@�d����|�� [l�T;���|^^�+}T�{Y=мJ��x��]V=�IS��7D������o{_le�@x�0<<�e�R
@��Ʀ��I�Z��W4'Vc{Jq�Ukg��ʀ=?%e0W�-�TT=�	�!�fy{o�-+#*�S�OH�)� k�F�,ѽ3�L}k���n���G_�,}^]�Ԉ{|������yο-*7����U�j~�afh\��^"��h�!�`؟�l��?�g�MMc�|�S���X{7�E��!�����r�~��ۜa_�}�p��&��D��%q:��~Wh���05����v�7��Qskk�
Qf㦡!�og�%�Β��V��t� ^�kp���v73�E$��F-v^�.�*r��NbX�z���>r��y�5���+�9���9�֫Ƣ�z�x��]�@��E�]���z=�N����%~�.��"h)+�ѿ���k�7�W�u�����e�⹠�1�}�?��V�v�@g�Y�a������%���כZ���a{?pt�n�3�j2\>�e(oí��8�*��e��CU�sf&�����3�R�o�^=���ǡ�^1Q:V�n�z'B]�4"Z�\5�zH\ݭ�1�q\7�2�H�}������������O������a�	k��\�1������ȷ'<��S��VئҵJ���`��lu�f���tAK�a*d�$����f����V�8�zK֓�z�V_C��kj�g�^�l�A0e7��F�e(�͝�ga�5��i��ʘWk��zT0�MH�	p�۴�f�Fƭ�EFF�W�4�z7�P2[��`st�c��:S�@C$R|z��X��#OG^%�/)�vr��i�	>�v0ʓ}��S�U�+�Nf��V?���[�M�RG�;�]��m�mG������2��;��pk-ǳM>`���`'��X��wTtB���X�g�/�+�4��Ȓҋg�c�Yh���.��7Q�0?���U�S�zw9W��C%�6�u�mƵb�0�+Y����������
H�h2����*u���Y�>(iS�(�ɷ����4B��u�Z+��0�����t)� � ]�I�	KoL
�l�y����)���L�whm��<��-��>��=z�$��"[#b'��9!��r�������OO�h��u��vuᑑ~_��i�����D�~CNS�z�흟J؍�Pfa�~�ϊ�xUk�2�K�� K�U5�B5t�F��z�ќ�l�zO���w.�{�oj��1�xlb>3��b��F�4˸�i�D���k7��UT�X6=Dv�O�Z�2��LJ�94, n��P���L �}���mu�����d�o�K ��p�s+�`�z�gup��,ڒ�J����o�)��6��u��dw6��m
�gf?���o���<M7(p,�b7�碨��_��נ��{�)�d��2y��z�ɛ�-�2�1�g�72�"�r����k/��g���hA6�.*����T��IA{�P�4|>i���7=�%^��0d����J՞+����y�:j�I�h8w�OT�n���^�^N�s|\CZ�劻�Kp�zY�3Q�):��źC݁
��ƌ 42ji�*�}S�!�"����0V-ӧ;��e���:k����U�d�w��[\ȯ��dzzz�>���e������ Ґ#	�Z��N>�����R:C������@����ki�����e���j��1�F��\���?�J�<Q{�rO�����B�1^'m�����A�d�X)9qc��ai�w�j�gN�隄�>s
�\����24������5:��(Ǌ���d-�ޓ�=���rT�,@,d��FU��E!:S~���5|c^�-;-���:���X�)�4�M���*�0J4��n��Pa��o���\��g��ե+�z�[�)�o����Aw�f�KpK3���蘏�<���Fi���O����3�ҝp����,`-V��͊�5���EQ�n���y�!Rey)�ҵ���վ��9��j��*��v���j�Ǒ�����`���=�&��h����8��-b6m<�I��nq��9��Zb��B%��[��n^��l�%�W�۶��O�����)���pa����M\̞A_ix�쑋 џ���^�!��&''g!��x���">�V/���1�__��-H>���`l�;!}0\��Ee}ˋ�n�y��:f˻�j�)��� x5�K����u�pu�F*;p����%�@p���Hj�W�Q\����W=��������X�����Uݒ���J����G��ٮ��J��� ���DB�ʾ�����4ܡ/���%$s��5�N�fj�m��$�_RYu-�*3�gdd�J��l܋�fz��ʪ[��'d�U5;��td�_��?��ų��i4���� /5~��&b�.e�"r��R�2�Ƅ�A��FE]��%2δ����7+�,)�<��N���։]�ϯ3"�u�R��y�<����h���g��A�hr�ʡ�A�W9(�&D&��7���L�Z��$Ξ�o%C)�`0Sg��L��m�g��u�`W�ISc��W�|Lc4?!�4�ֶ�R��$U-=�N����g�r]�B��pq�ʒ�32d((0��B �{�,l%N���F��s�Cw����_G��^ʰW���ǜ������tsSl��͖�ҹ�q��W_=�[�	F<���N�5�Fc#�A:�J��ҩ�%HP_O_����X�����Ș�[&����y�n�-A��C����6���w�(y����N�a[�<i6��w(��q���Ige� l�4n���I���V�Phfӎ��8�tw*)�����Mӯ]y��Ap���*���#�������4��bq���snE��u	\�V�i�/PK   ���X#X;Y�  �  /   images/2d4ebd0a-2d28-4b22-8d08-8a7e71760a75.png�XgTS]�N.	A$�

HB�N(" C�.Ez��BhB@��6���4E)R��@�b� J��^���~�f���_3w����9{������y�jaf��<���`�'�,a0�$����9��xYꧫkqRWmL��;��^���f}�iz��J�m�&=����a?Y�}v/� <t���=Jt�O�I�=?#�(���|;�3�,>5�>zT'�ǈ��y���'ECy�xx�aX�c�����'�0{��O��
��)��a���{����z?{ۮ��L���<7�緥������$Q��\���~�JL:1�fa��~!�7�c�O�Ud�7{�'�|��J�,;��H1 �k��8G�9V=tU�s3�� Is��at���o�n��mx�y��Z�i�%�ǆ�R�Xߎ�v��.��%.�X9c�c�1s��[�
a~4A���]��πcʑ����B	s��ꩼ��� ���Bޛ/#�x�}z��nֻ,�T"�LL�������џjV���Ԯ:Q��Y��v<�%�B0�s\J�њk����X\�qgǝ2
����&i7{[��k��~�p���p?�S��n
eB���'�p��|�@]:��?%���⎠v������33��%�
�ʛcW�vd���K���޷���S`<n;�m���k%���!�q�Z�0o�0"?�V|���w�Z�4lE:�V�V����`Қ|�ΪO���}�\���0
���׎�S��~�oK��y�v��;��h��W'�`�xP��=���n��O2�ˍ'-�� �.����nA�>�+Nh�V.d�}*��!I���>�f����q]�{���j�8u���ɱ'���8���i��u@ꕮAA5��]��o�(Vs7�q�+⚩�䁛JF^	�d=�Y��#�_��ﾑŭG��OX.�"���Z�K���{2nI�ʽ��#�N��9�Hl�m�vH/�^�{+��d��7-zC�E��Y<��0�(`SN^%5{�z�`w�X�(2'��2#I��O���}��9HpOa�r��0(贫V��;�;�M5y=1�չ�%3y+�u(��OC���Aʰ�+�!�D��V�>A��9ƹ�;E�5=���{U�j~S���,�lnrrrj�e��d��e�����S��D1L�����_TH���ԍ��wgX�Գ�j��b\����o�n+��(�j��nm�-���Mq��_?Zo��^�_6�CН7G[�n`3��H/şzj��0<���EQ���w�/�y��꽭f1�>(1�>�2k��o~�G�����d8�i�M�O����"/�%uK&���������[7nU�P��l���pOx̫۬�S�Y���
^�JY�Y�:�Zld�haj�x���g����+&��_����8^rp��9���N���:����]�U����c݇�̇�[dL�LU����|G*$���_����n���a�GJJ'K�>�ҧ>�u+v�w���Gw珷��������8������"՜^8.��S�$*|>O?���ȣ��{�b�3zG�U�����IV)�8 ����|�˺��M)�t҄��ͤ��}��,���n}%�,��;��29�wF��it)�R���h��h��A���^����gu�ˣ�B���Ǵr��q~���;�B/��1N��RپT�[����?�ۥ�r�1Z8׈�!!�5��V�Q�6:��C��ه�3o��ff�ƻ3g2����T�U㪦;y8]
=����t�Bׅ�BA;�ŔR]j��1:���S"���M�؜�b^r�8�x������O�񊖢������ڴ�W?��}��-��E��\�ҍj����Y����#��v{�O�	�O���i,�,]@��]��n�iqT����B܋+F>�\E���Zp�:�%V,�$A4]�e�y���F���:{*��O_�P�Bs��Pے��K@m�[�4��>{��2k�;us�/m��z((r+V(����ue5�b&�3�1ڢ߅O�L��]m��j�혭2�u�5�qaϊUz��7ݤ{��$�������,g��|�^�}�e��]�����H�ϬJ	�	��=�e���țS�M�s�g�ğk������-����r��c9e��s�Ů���9[�pϩA���I�5�/��_�4Z&�?Xq/R4��c���\�|?!�s����FLS�lzy���5:'���ڡ����R�^�%��ӭ2u�Μ��\�	O����t?����t2��k�6��b2~�<����VH���.ma�`��L�W�F^5}w����z=K����������������׹7�mɭK���M��t+���}]J�ލϮ�m>��Y��_T��y�d�I*�y�G�e������c�c2*K**c}��N2��~��"����ZH���խ���� �g�����{�~{�w��,�Z�M��`Ϸ����׬��Q�4[wZ�ȟ�â�#�Y5Y!Au6�kc���*m���.��L#�Z�zEQ�-6\ᘼKHC�T���sU�jv�W������E�e>55	_�6L��_<��Q.��b�G�EO{w~̛�ڿ��#�e�n+c���fk��j���^��K3�{t��F�JU��<��UG!�\xO��������>#>�y���R�
,
�oz|��=�~�2�Ŋ����
�Cן���_IYi��+���&�7�kn��r��o�����1�c�VgWWGư��|ה�ʨ��%_i��FM�!�����a�4 �
��`C�_�D�S�lÕ�-����m�4`��*:�q�Cr*�k���:<	��~_���{��Pܼ4�\���]i����gbP�v�f�d��'�>�$/��ަ�0iHF�@�A+$�����#��%a,�e ���7�������ӳ\O��AԈT�_��*�?��3m+ݓ'���3��+ ė�伲�ڇ�`��w����d��gmjgjr̓�/�~���%O���_�x��B��D��!ǈZ"�5�A��0V�[%������Z��>*� � �C��h��3��,���6��D|CC�a��������`����:VA	��$iȅD���BD�,�u��B<��C��{wP-��u�\y���) ��mA���`���������1?��y{=?(f�����&����o-��=����-��gK��`]�?4��w��6�ϓ�
��D�O��������3�V�FA?=sk��.+7�I��C�\��3N�i[�� �{�f��4<�*�E�P�(����k�j�w@������������A<N��ÕZ�=Ze.�I�ZΛ���kEo�W:���{��I08 �����Q��Qh<��'O	�w&b(�=�+$��hz4׎���+T�k�f�{>��J��ߏH�����ZO�]��p�Nii���e\��F6��R�B��Vӎd�S����]]����(=*��`۾;��Be;���HF[��J�(�Eɺ�Y���иLbAFl
�������y�x�	 q����2Ἲ^��� ��G>��Sh>�{�2]����4��ho+bGeqK����w�����,�M��ܞ��Nl�e:S�*k��m�~��.k�q���;��P��h���C^�l~(���:�[h����͂|p�_GxA ���P+C�/O/<�ľ[��v��t-�g��s!@�QL�DB	��:L8��T������J��� �w芌�n��Y��d\�?��5�8�b��Jb�<���g�G��y�t�܋���eZq���x%1S�#~���KȌG\e�������݋������R6Bg���X%��p̡@I#���W��O9�Ye�OgL���|�.�G����T}��0�)�8�����<E���
�ɛ�q�y��E���Y���Q]1A$Z0��i1LXG��
PƵ����������?؏����B���h��1O�3���m��L�ע�x0nE��mq�������M���WC
�LT�����M��8��+<���tSN(�����N�PW�f�Gւ:�k�yZ��EQ����@ 愞�ݤe���9#&ּ�Q��:�#/��Ր��ul�j���8�
�Ư���ɗ�&��ۄ)f�>��/����I7p�FQ�,��*����#j�͙9������NĠ�����ƭl��ku���hz���_�F���[�J]�b�%7�=QaAӹ>�(A��㲦?n���(�Z���_o����_�<69m0&�!,���"���``S��/M��qP,&�������������2:S�o��_������|�ȅ)��9��R���l[sȥM@t��O�>��x�>��g���E1��#l|��[Dpm�g��7�|�yZY��V�=����*
� �A]��_+;.�U����Z� ���I��/��L�h���Ԩ�Yd� ���x���JgN�D�>;W��E7@k)꣭DkW��ev���ˌ~/esKG�GM�5>qYՎ�?𾦸:�(�0ч@%JX��Y�^�fG,4��q�Pi�'�?���;Ҁ.3�{fQGs�n���$TcS��U��b�)b�?Ă�����Ǣc�b�j|`�mJ���j|���!V@�������˳_���(sj�q�D�baC9�ם3ӟܭfst������`%�oҘլ����cd�H������;��{ƅV���"<�.�qD���zڡ���Bs3����/\����<LXGV��oG Z�Ʉ	�ā��k�1��D��Ṏ��B�i�v����W]�"�:�65�u6���N(�#E���խv[����TzZ���O��x����F.0b��ْspL�����X��T�����VX��ӛ$��Qo��j{L�Մ�"݈��`�ȹ�e�QJ|��>��ݶ�\���kgF���Ix�/!��3�y��<�NPEn#�]�C�HZ��n��{u�V>�7�H��5�&�r����ț���G���}(����k�Ʒ����yCt������Z����2�d�����}��Z���x�������� p��3ᥱ=����~w�Y;g7���{Zˋ=�B��p��D��o���u�� Έ����}q�w�<E�,g��� ��(�ޕl)���
�$�p�Z�����D�������2��@�d{�������r2��=�w�[�jb�
�y��so�V����.�1�Nq1�4Y;�O	)o�*�Q���)k�-R��p.k��������K/��︂�(#�6�4�;vD(�[D@G*ˑ{���˻�p�<������W�ȧ1]����G�#C��7>��|��%� �Q�㏙#��c��V?-vR�n��S	�A�0�����n4��m�^7�������s��4S���D��M���1�ʎ�����_���^v_xZ�G�Oe��ͯߛ�ƁMd�웁4¡%pM����l�fC��5v^�����2�N�nK�ԋ��v֕	a6/�y�y��}kz����l�`��ňvg˾o n{���x ��rQ�}&m?y�ő�<���g�/gL��1�	E�cZ%E~q�xm��Г:��K�t�v�m.`��9�iO���AȢ�XT?u� 8g�FX#m!L�C��B�T�����#o��!n�E׳B`�$�?����BPs��o$��2&�ӳ 0,v�+7���b��Q�|�2�1s�R�^@��+�u;�(������\7���>^~<u�l��K �F�'(�B�;���!L��s�"!`b5� �B�
k��Շ��j�wH ���$�Bo�J�#g_��:j��r�Y��_�b^MҔl9pgK1�q��n����!u�g��.r��fE��1K�f���\1S�w`����\���@}��V��U|'��* �"��g�3��ͣ[��W��53���XM?f*�ȇ����Դ�n����zO�KI�����s#���R�D��z��0��SH�f�.yM�޸Pq�u�� �����_ns-,���
���u�m���XG��Yľ ���&D&��=U�FQӕf��O5'|�g�L4؊u�T"~@�t^9to�"�R�b�@�0/���s�*��sw�������j.� b7�V�/���k�&'�R�j�B��U&��q�w\�=�}�g֚��j�1�ߜN��A�Ņ�*���N�\]�d\�Z���*<::�4���9��F���
�m��8o�OO8J�5<�FL�G1kS�~�KBa���.�}��Q�Pm�O=*����/o��x�es�Z���Wi`��E�v���Hra�aQn_)~O0��%D� �&n7H1>Q;u6ƃ���K�ԓfo{CGӿj���Ȧ��,M2�u�11���ضW��b���.�gE�6����.�Ӏ"�%&M�d�ne��Xv�l�Aizߘ�|r/��B����V}�*x�ȴ���2��&U]�Uo�}�u6�,�My���xUIs��%���VfX�`�d<�)� �+�n��P�zg��!z5�7u�bK�i{ ��"I{�sRfǢ)F���jdݱ�R�P9~�o(���
	5M�?�C>D��i����V��Ll�����)���*/U���Tp"�������Q�VX7��6�7n%={��~.��x�>fIx u�u����Ɖ�9`���~ێ�_P`�{K���Ӄ��B�2kˇ�fԧP:w:�F>�0���]���u,�Եf��L5`q��F��+��&���
@o��|�R�;�_�8�i|���Y0�a���H�e�����̿�P���u�xc�(E�Ai�����v�ġ"g���ְhn�ϣ ��W���f#��*�(D�X4��1J4Y2^ PjE�<*m�
'�����+ˌ��{Q�"�!})-��O����`p���FM��J��[�t�ź���t܊��e��^6��K�!?���+L+����/8�	T��X3�ɯ'o��\�%}T.�[�~��\{���e���"���V���댧V�k/����|��WغOk��^c\���jr�^��[� PK   ���Xt�ʰ
 � /   images/3243dbfc-afd9-4800-9031-ef944cd75f6d.png &@ٿ�PNG

   IHDR  m   �   ��l   sRGB ���    IDATx^���$U�=�*WǛ��f��C���H6#��}��>y&T�
"AT����i�a�o�����>����{��'ӷo��S笽��k�֖������[�?|�}8E��AF� ������ñy3p�{�D�E���y���Q x쑍���;1�ː���:�����s���O?7�J}W_}��������[4D�	�	:��1P��k���cӖ~:";A!���g �F��srpu~=��yD�MӐh�� A qF� 	}���|�K���T���^��.`j��� h�#\~������5���=���.z������T��t��݆[ޔ��p.��쵤����q����w����3O�W�X����]ԡ'���~��c/<��F��S�U��-�G&����ِ��� FOg�&+�~!7���#�kH|5�zXB3�@��QY7�t�1uDq[K`�:���g���P�d!�B�	-j�2�i��9؆�D7�tו�l�@��<mmyLM�D	2���YC�5`��(�m���d]Ĝp Q�usp�C�{�6|xA(��p3�Y^r4$Q�|΅�9b ��LN��^�J���64⚼�u�V,��M?Dw[7���	4X�� 
�5$�-�kQ�Πֈ�[6&&�(�30-�f����ӈ�	b������M��p�,b�@3Pk?}xQM���\�1�i��I��KB��������;�4�鹍�E���`#B����,I�!�Ԛ��Q���7H��Z�J�]W�m64��C�~B��z�`(��	˨#�<qf���gP�P�t�E:.��4���chK��/�Yob���Ѝ"�}r�G�t��zm;"�-Y'� Lǚ\�$�z��H�v:'�� �L�|u-�f��!�X�B�$�G<�܀��C�l4=A�A�-�Ն�δc��K��iXA	F2�Fi+��(�DCir'
���Q�5W���K�w�<�l����.ڲhk�%�粋��a�xӁ�jv���8��W|59�ؾc3n��UpR���Oc���ӛ�Al �a=0w>�_=��n�'2�&�<�|�Ñw	�&N:�k����r����Y�����Jx�5�����!z�:��g������m#D�L�����c;�H1�������k��L���0b������U9v�H	Z�,�0G$��6�u$�=���+h��Qo�?�����|�L@K�(Q�;nt0k!p����9�h.�����O��_y��ˋ��G��K��Dh4�x&~t�������ão���������߅}�Z�#V�V�`X2�Q6�]w��ig�FG=���[���Yq���ь���v �.��h�m�,��Dq���ux�ڠ�Lۆe�Rԓa��\6��*��f����	#�!1�s\�A�����%��f�\��W+��78�Y|�N@�4�� &
K����eY�{r��mC�;8�0R7h@�RbL��`�YX�����>
�G�Π����C7,^J�4M������ζ<�(��5/��5��s�|��J�Q$����]mbhB����HtIl ����*�@�7��e���b-[m$��"M��ƍ�{�#t�ӴF1B��</�k��,���(����;�4�\I� �xF�8�[�O`bDI �4���ćf� �"$f�8�q�ah:L���!�5~���g��A7�6@^�~D�lޮ�M��>�\$��kh�(y����☣�ࢳ �TԠ�l]W��1Ĩ`��x�o;��9�0�����D�={�D�]=�a�������װM4c���h�u����Ԑwۡ��8D�ِgmۆ8����]֩�0���^uh�|V� l 2�>��p��A͛u�A ��V~ޱ�LVc��\!������u�'�������1����0,]Xh�c�����-���D#,�R!�bh~���x����2�W�Z�w�������W݈4�\꘥K?��^?��G�|�<DMܳm���Mm����kh�:��O�'�|�0�6�X�'Nסr̾{-Ŭނ�������s<��k8�]�{<�$Je��B�ǉg����w��,.8�8\뽘�(@������C���u���aG�����1$ZC~��gO��g,�������oA.���>�\r�p�߆e@��r6�ۊ��.���8����+�!JL�Y[�s|���vxq������7�����O~�#e���C����)�����������'LT=l޹탋���k��?�r�kh�F1g`��v�^����YzVӰ��^�G��o`OL�����0MQ�A-��/�I��Z�㻲&�8�Y�^�Q�8��Q�ë4Q���������^�O:�vnUט� cm=�h�A�q`$�l����&�l[���`tb
�e�uvvt��y�ʄ����,7���wgP�ֱc�6��#��[��� �4� ����ӣ �׽�'^}QW=��l_��b[�� �r�0SxHw�>7�6��{M��M �)�A�@J�W ��X�4<�	�K3��DC�Ѝ�"It�K��ȗ��7�m914��nh`h.�5�KA��Hq�_�p�"����!�9>����7p^5?��`��\�k�T�>���zV�V'��(�O���q�1s�,��]e�1PT�����̞�.o}���T�`��=��	/@��2V�)���7�;:Q�V�Ĺ1F��~Z�L�1s�q��G�g�������F	�ԣе�n����n9h�%��hK�7���zZ� ,>��-ؾ�%8����9�/F�R��y�c�N���5�p�Q�=��_\�y��������������x����31ᷡ�m`(l'J�4��K���������-���1��/<B~��!��w��������X�����X����z�����C�j@3m��v�����n�a�p�ɗ��}w8y�w�8x�;?x
,x��M���W����~��::��Po4�O~�������p� 7��VL�(Ü��rţִ�,V���Ą�G��
�j��{�^X���>_xk_�ҵ���Ħ�[q��.Ƕ�[q��{���C_�-��D�T�5?��=j	L���7pӯ���hk��=��o��x��L���ø�w����dn;vlڎ9�z�b�����wwb�4�����o^\3�L��.���7o�{�<[�oƃ?�\jm�:a�w@�����܆�<������c0�. �õr��5��j�m4*%T�ӨVJ���B�@��tv��Qe��h"�|�~ ײ��p!G���B��o�ycC���i��w
�t`[&�J�e�KX����9/�W^ZõaXf ��b���c�6E�)�2�����W^�ߍ��#�@ej
��0��f|�;�B�|����vy}�G��C�S�q��z��lQy�j�����l�`DaӠ[�2>1ʵi�Y��π6#	9a3����&�	B=A�Ώ����kf�@��!b��<�m�R�4���#��	܉_zٞـf(N��3$�i8����	)�$����1t�/�C��,y?�G�LG>7��t�c�� ��A�+!��X���.8V>�eQ��Ğ�zA��}�8����U�|
?���2F].ۆn�`e\�k�@'&�@�=�HaÒ�K"ME0�-bz�|�\��B�8B�B�&@3`��<l'�#>��������H��[����vnx��/n��!|�C�a��8����lkC�R��M���P�+��hxֽ�F�T���Ksp�w���K<쉎��a��@����$���u�(�s�%�|=�{`tr;n�ӷ�h�\lܸ{�3��:N?�c0�<�>��!�|�<�����k_�^-�8'�a�k�+�x?��=���C�<�_��>�0�����j��D,�݋c�_�J	��g��5on��`�y̛5Wλu�v:��!~��"����S��_���Q婗L=}]h��F	�tq�7ԧ�1Y��i��C��O�RT��~�{�s����I'���;	G��0�S���?��WWmEww�|�QX� *�g� ��0B^2�%�)���_�vnņ�i|��7�{mv����wo�y瞁3Nޗ�6l��?�U9fה�%{����%��\|�g���<��0�tŏ������qk�gV�ř�Z������op̑G��h⮻C�5`:tuϒ0ܲm��*:���D�^C�r�,��!�u�r���Gbx���(�`�&��ctr
�6o�α1�b8}�r�[ �q��ɉi��u�^ C7��8&�'�l�144* �7؋=/���3o6�f�Z�f6��:Y�Y��3�oن�{�l��\�|6�,���Zc�2��,lS:#	=�z�%<�������9s�̆�wa:6l�в144<�S�M"�K.Uq<�D<�8<�
X���M�\3ⲴrD�.Q�
�T� �h�6�X�S��DG����yO�S(E�p�ӧq����W��}l��ЁfűI4����!�Xy��e��h�:�#�EoB����5��c�}��~`!!��+0���)P��؎���7�w�z4v�ǁ+ Fc�j�r��o�ufa���yd#��ö�mp�@�bpJ��#�Yo�k^S�#64�M/��ϑ������K����/�oZ�Z�Z�0�POs+0m,���Sص�E,����@O[���n|�s�M�5	���i2�"�⃌�=�8��s�F�X����k��O��;�{���:��:���$�����V��.d�Xf�n`�<�cO<߹��j��G_���^��뾍C�+�	G}\���t�zXsp���cǸ�'w㟏>�f���P'
itT�v�?|��a9.n���������q��N;+W.����=�.��9x�;Wb���l،������ߋ;��2��I9�37���W�'0"�Oz����|�s'��@3(ö�X�j3�x�#x��Mh$j��q�a��>��	�����z�wc�!���|;p��c����TU���3��������>}j�x�%�����Ӻ0������A��ء �3?��S$.����j8��Cp�9��x��a�o?�m Ԁ��l�t�!��ʇ�o�y�Eh��ފa#��ӰPm�l��o�^)c�e�&joS��V, �ɠ�Pm�{
K�o��׫�j�:�iy�^��Y=�׏΁�:P�7P������ �2s٬J8���^4|�/I���y���_+T�,�ïB��")�d|����p���ƞK����֚a��1���n��ӓc���{a:mX�h���`�\�,B[G�P���$%I�$��@� �!��?f�6l�4�7�aJ�P6#=NrkҔ�fR���A��=L�Ͱ��͠�g!�thq�K��+`%��ܫ.��mu�[��}#Dd0}�J�v�<Ϙ�@�!d���Gn�ϡ��s��R&I-[��H���~h#�$��I�2F�ZE�{汋p���렪��]��ǁo_s+ֽ1�B~�{���j��:a�a�M���ȕ�&+��.���|f�r4���L�YK"�t*�K�[Ѻq!�i�q��8��b�����Q��ߑys�U|�C��5W��f�O��6�%��~�T�_-D`��E��<�`p^�HED~X����3$�����ȶ�c�T�M��v�H��������`	u���}�\�r���t�~m�\�3��z
�^tu����J�O�^܄z�C��q�9����A�-[W�yt����R�'h7�/��N��g��\���w^��ɺpl�f��c��i'�d��~�fw�����E'��q��>��p���q_���D�`Zׅ���4��F����0��ڑ8��~�Z�������O`�hV�#��	8������z��v~�99��Q��'u�˟��>�F܆U{��#��3W�1���w?����(eL-�����g��|���$�:6	�Z�>��������{�@3�X:7�>u�����U��~��x�e*1J��������/DG{q�]GYK��ò薉q�e�{�Q,���9�(��h�I����Qo"c����e!N��9�f����iIf�t!�P-���.8n:yY����0�[��(
C7P��P+UP�)��{,B��h
&>��&T��ɹ�3�����k1<<�����B��;:���9�&�Mm���0�M%���A�T���`n���f�1�:b�/���H��֠GI�O���f�A�-�fp94nz�As/� f����R��91R��b��gHg<m�����-�6ȗ�M�k��VÓ�%B��T��w�Z��M���St/��i����qs���Kh����=�K>t��k6�,�����/�g�7E��߅��c#��VJ����lq`B7����E���A3w��"4u&bi�8�)�-D�	���*z�	<bXU�2]���,JMޜ��Z]�=��Ꙛv��h5�^ԍ��!\z�����Ȁ-����P�O��\���*����-KI��ި�W^ǃ�<�#_�g�*��.����&��D�ni�����bۦ4�@&��9���}�D	�ׯUV����k[q��?������<�CJP�lB�g �=u��43��$O�}��a����t�_���~y˵�M���~��n�B"=�! v�a�k_:����a;tO�v��4_xf'V����i�O�5���k����٫x� �P�\Kwa<41�k��Nh������G�����;p�]������&8��{b��S��O��,��ٻ���M��@�$��e'b��	~���?�W�n��q�yC��៫ hֿ�<�GW
�_��2̨r����	8�݇��X���g�~E���f�F�k��g�T+eԟ�1/ß�9��&����8��+��w��K.����c��V྇�Zz��H�'Ȅ%a���:�S�S�(t�tM�(�kGG[I#��	GZ�5����p�A#��8��3��*�ٷ�G���U�Ӭ{�U�r��$~2Yu=�j�
Ƕ�7�m���qn�2Ѩ5P-+O?aXA�a�B�j�KX�x1�ڋ�M���M��>����52!ɥJ�7c���'hc|�6��]��P'�������"�[�3x�T��P6�W��T ,��Ꚉ���\pɅ�4��߽�4Vt�-)Z&�i������m?&Q"@��NEż5Z .�K��)B�"uc&�p��E����k-����g.����"��糩N��C�>�������Q(	b�5�b����s��"�1�U�_�|:���ۛ�{����qk����&�vu�mI`��tO@[K��&!BF+-�"T��ٝ�3�D��y��*<cָ�ɍE�?��sv햇�V�9C#kq�����=?�`G:,���՘W�U"9T.�.�T
�(]�9׌��<�J�G3���?�H��y0s����k���[�+/?��ތ�>�79`�X�☼^�xn�E�|X�p�;.��ŋ�|�}@�\���7�|;G��ϾGtӗ�S�^����N��)�>u�_X4��y{����Ÿ�>V���o�)(T6����O�kV��_���'�����K���7�l�����;����<��"]Z<Â]���K�L3Gs�u<���x��	,_�%��M`����@Ǒ��|퇧bő=(:e����k�skG�?�{l�����92R�C�?�_��ohFe��6��zY�k6Nbh�(���=��4Q��� ��{߼��P�?�x5�c�n��<�@>�̜�	���U�c*�R:���Eo���f"\�'���¨*km��%���Л$��Jr�� vr��t�F��Nݻ�Z�1�1�C�V�,�eS��%1�=�4�9X��k�i�8    IDAT�	��f���7��1]����=�9tuv��y(OUd�SQ�$���p�ٜ�f��"�.ִ�:9h���m�!�'ȴ3z���%�H�2�n��(G�y|�Ķ��������#`�$�f���jU�g��j��%a�j�e�(�UT������Ԭ;��d�1�!LUOr�⬧��zCl��is>�-�?�ϊ`�Ħ�ί<�z�$Zd�����!-ĤO�c���&e@k��ǺIy�Z'-���6,���S"��ITJ#��%'��C�V�w��>������LB�~cN9� d�XUxM��{*�������/"�4����Nm���FX�9h���$T�Ċ~�0i��?�fKW��+�;����V2�� $=fpmN�c�0���,\6�����3�����XZ��+Cs�ե!��C�X$��Օ�w$���b/�A3IF�شy�S�O[X�Յ��+�M>����S vm�o�c��.<xﳸ�_@1o��GY"��>�Sl޴�I���'qҩ
h���m]�a>z�Wp�I����.�cXBI����q��%!��W!�oUq˯��׃s!��m�n��#p,Z�����3�k[�����S��'������G�ſ^��tIy�:2�W�<.����(�D�#
zc��
}�K�1��w����߇�	\����W����$:�;Q.7^�8�e�~{����0���;w���>{�O|�G��]��W��}��5������X��~��DM����߼�"=��f|�+ݫٽ��69�lf��*�^��K�0a�1�LQjݽfNQ%A#��ހ����4̀P���xLnp�9���"��s�{�����t	I�V%j�ná�5��(��Ӥ���u�� ��7C������y��K�q#X
�eh	::��/�k�Wj��
LR]�*�<�9e�ח���w� bh�	����:<&�5���+�-�h�F@O[Q<x�0��( �l@�3I�#�ȽHh!J�и���Q"0'��%\�s&n��CE/�P1�0A&-f�kW���%�.T]ӌ�:�L�򌇝zڜ3�
�j�H86�h�OX]Tb�~F&�h8(A$h3��s��N#z�⫆6�F����4�?���~c;�Y2K�r�+0�i�����h��e�p���kk����h/vCk��%��hN�~y.-��ш��!^��:��%��)���'\������b�ԑ �Y�5��5��
[W��@v�u��TDГ�`j��I���GDC��DQ ݡ"��Ч�a�Y�`�y��IX�2.�W�=��X�c/P�1��7�Ж�����ꯞ��	�}q
��X����ܪ�u�6���'/�>&G=��į��=��%U ���?Jy��w�M�o:3��?��n��q��b/B՛D->����퍨	l����q���>$�To��J��ûNP�������W|�v�,�c����ܠ=]���LM%�B6��]	�Tsˍ�K�@G���c��q�G�Ǔ���1�)�H�����7p���?Uɶ�܈��]������s���;:���|�s��[_�{,��~��|�T1q����00P���$U4c��q�ʥx߅�b�%���%?«�G ��lC�w6�T��np� ^��Z��l�T��pmq�i�R�ReE�G&`=��]���nZ}����&3��h(�Q*����`��K�J��(F�5%���
�m�p"�1=Y�t����khR!)�g	��P,fe7��gEd��"�S�j�kzb4��6-t�)��l&F�F��ȣg����(���dW��ZSk���BZg�����C6� h����h�v;$�H6�U-��
 8�\o�� VIr0!I/U<�ԳW:�gPQՏ�:2���T��3&}A�$5�6�O���zt�w'G� Zq���+/]�N����V(@�L�x˰$�khQ C�lZ:�Р\0���Ԉ�Yhб�tt'�����|���z.W�b�a^�k���z6�����o}K	ʍ4#��fs3��a�#�o�-�"Yԑtdy�[s� �		V�Jd"�L)���)S���>5�r.���[%|��k�+hhsIu�0�||L4�*��ȳ
��)z�	J�U�hB;
#���*��C]s�J�>^~��5��w�L�����U����Ɍtӽ�PЌ�z�ɍ��O~�U/nGߠ����{�
;wMcϽڥrM�PLH��{���k�Ǔ���Y(erB�+%LMN���7ޠ�]����s�`՛[���F،�]� �YF�7{��я\����`���k0��H���; ��5}tw�	�D�$�r.�j�:Q�@��Ͻ���#�d�T@�ز~3-����&1�k� ί���]Y��߇E��v;�	�j#�A�ez��v�1�t��h�Эӕ��*f�׻���u娇>��a�;�J�qZ�0�� ����h�� ��!㺨�j
����v$jf�@���H��mݑ*97�V�%�a��7� @<���Ra1���`&y��a��d�
�<��'BOp0;��8�0066�Z������7pM�˧��ؖ��8���ec�M��Cc��&�ГD���<�:�܋r��zcS��pP�R/)��8�l[V��|Gn&UA�v��JCdY�,�$Ʌ*&�l�l#�$֨�`Ţⵉ+�^x_- �:&-�iy���hI�Z�*�h�TO�,-�<]j)'+�Mc�;��Y�[������Jz��+�25��X8onpV�F-�`ٍ$\�Ȫ2y��Z*�4������2�-X��)<���0�_�Xh�n{)Y�ׯ�%����;���j�^D6_D��RF6�J�*��$ɪkb5'�|c���c�D�DDJbY�z��PCI{�4)9eF:A"�!�u��|�\��o}�DdS�x�]�
a09�r������)��G�h$1/	��h(���4\3j�Ke`#��o�cЖ�ݤ#[ǥ8�ϟ��UAŖ]�B]�y<���x�2�v����hT�`\��adrЭ˖�¥:���'�r��㎻��%��^���o����h8y$�#e��9�&~�����Ǟx'��'|�5���?Pm��f�N���چ�a���ᓗ��_t0�l.��f�+5�/����"rY��5%y^�!E�$#o��э��|��qÍ��}X�&���h��_��u?~	+ʚXfbT�L����A>�k �,�G�=K���h~n��c�����ꉊj������[�S<�\������cS	2�J=狰3.
��D.���4+ �ʧ�(%�>�D3H���_�=8h]c)�wsi_�t�/Kg��vuE��fh��ˢ��WEK�a&��&������ Ic��Ղ����f5���,��F���khogIt�ٳ��J�͛�K�"���t��JUf!���̌K%K��.�ݽ��hzM����f�^��(�* F��A���BF$��e��Rl��䡱��>�O�ɏ-hRXCI�;�F�Cy�,m7,�'&u�ۤ��=JQ�$��TQ��o�(@���3�*Sf�ru��[aj��h�V�οv�[
�F��{��CU�FN�p�#1$�+��v�5��&A��a^b]J�Y����{�C�=�>�N>�P|��+���|������혽�<Tj��{�Cc:�����֞�t��L�=Mɿ��ɓd�9E%�$m�8�|����VH],0���~f�?�z�*U�{
Ⱥ�y�F7b^�����0,�SIJی�@ �S*N�6��hB�+��Xi��"xj$�Wj L���Q�]�#�F'����l_%hp�-��oĢ�=��&N=�H�~}z��1o�A�~�s��{��g>�=�U3�v�8�Z�z[ԇ��/<�=�
���{��o�"�����UH�e���pq�ʅ�
�:�H�����/�w��̝3�m�e$�:^��#S�W�É ��g��$6�|b�\�Y^�l/�H(��V����MI4H��VR�ק�7����/�~}�RAfF��O|��R�]�PV��Qy}���p��+����G.�3O���Y�����=w�-�Z%��V��0�!v3Ȼ䷶�9�~�1������?�֬ن�����=#}<X R(��7udMS�j]��X��-9�<xz�r��!7�	T�H��S9���U��.a�&�i��oC��)�ɛͦ�J��"xlC���ؖ� �011��Y�P�$mJI9G�T��D	�:��P7�:�3�`�o�P�cxx'�t��4A�T)�����e9�tU������ڵs�-B{'���E���Vje�MNc����.PDEGl �iä��-B[G���զ���Ȁ�f����!GSC���P%B�����8��I^�I,k�)���1ne�d襧������[�=C��_Ҿ���"�F8Zk�s��JD'�ŵ�&KSCOm8?@���.�Ũ:��Y�ȍ��/B�e� K��1��M1�fbxd'���ȻM�u��8p�^x���D�T�͝����#�?�Ï;���8ι�$<��&d��<��!�:T~x���t4�E^��*	������V��֜�[h�$?��?):�Գ�H���qa$��**J0��
'c��&�<`:�t�A�U��g�)cr��8U�`�z�4�����g56��5��z~~�a�^�t��������	m���K�R�y��06Z�PyK����oV��&@����n
Zm9�;&�msQ-�D�5��ݍ7�����Q��o��(vuc���0sy��
pHB�����Rq��U�8��"�ԜLʔ�8MV�G5(!��מ�ӗ���^��ƹ�g��T%"�L[�Z�t*�"����攇x��+C6*j�"���s�=O>�����{�x��7q�Q+���6H&�����(L'F�2B��<�<���1���m�My��G��^C�c�o.�l~=�K�+���uxUj5!�?�P��jJ�&���i1A��y��Jr�%e��^�*I�1$n%���U�@@�$�9�p��0J}���uu�;���c�n�\*�ViH�9X��i� A�2=9��;���%%��;?F9����p��+�e\�LD&������&����ӏ�btt�f�1vn� S)� FT�U�_w����w`�+F����f�x�ŵ���6�D&��>�k�˂��Y�;|�	�ɠ�/��ș
3R���.�O���ץ@���!hLα�R�nL������ �Cc9������i��gf�R)��[>������V7��{�B%��LR�+-� A��m��?��ƄFz�|='��^ljS��[�ZA�*Z�6�w��L�0���>��nV�!�3����5��+T�~��O��w�6%��"v�`�t'��$�NՎ�UD���{���!SeP
�L^GT=�\iI^���	�MߗA��`�c�	�[��a�]'�/�u,����6�֪p#�)R�oI�Ĉ+��8�T�¢�J��F)Tkl���}U����4z\�f/������	Q�MA7���78 �<�e"
�WD���Ϡ:�Dج�>��v�0�c�3κ�L�]���p3��R⤸g��t]��P�V��.�ti�՚Hl�Y���r]�keX)�s�lJ�6q���0�I�Y.Fr�l�ê$r�Lte�:|C5P�E1�
<N8ew<���&j�j�X� v܍��![d�4���(U&�grof���|��Y�155�ys�R����)��~�^���ieݮ� �b;Y��QD.�+ћe�:mmm��jL�1��n�K�+�J����h�x�$���͌8LTrP-��G�FKw�'�1���U9��踀6(��^g���@ܬabrL�����(�c�|9ǹ�%�{��Mb���v�3D
�,�߾}�^˖́c�8��C�J��֨ضmDz��8���LO)@ظi,Kþ���V���+����#�Ӆ��_��aM���Br���nۆɩI���vCWO�E�1Xk�D��,_�c�=��nJ�!���>w�@���T*"�>���TCϸYJM�-����o��3�ʋ���?��OlV�*���j:+��^?��CXqz��F�V�I�Jܔ{�:;�@ۆ)��$�$lP��m'ق��-]�4)z���������->=ń���:*�whRn���tF���ϫ���x,���ێ��ALNUG��X�u�8�z!w�V�k
ԺWƔ���Q����sY��H���4���C4|Oh.�Qp<Xz�}��2�nᐽ�����1Ml��O{��<��E�EJ�. �T�R\�U�oC3������?�K�[����2���]�r�.z�4�L�A�k�>�vm��9�����^Ε@m�T͈]�b��j�;��Sp�aOS�"eS�~ºhq54*>��7bg��7-�0��T����I��e:l ���mg[�r@umd[�ׂ�ht��d״V��
�P�^Cgӵ�%�ln��!�낞��M@�˰ru5D�M�	���(a��I4C�麀6��̚5W6�c%qF�ki7y-�f�)m�i������T	z5hN��M��0 )U�g��|�XS#��8�ʸ39�^��7b����)\���5�n܄�΢�w�>J�519���~�����I�f�(r4l�6#�����FF�1�}]QV���sO�c����B.��Ĉ'��JI�L�/9���W�������c��X���Z&V��ڊy��>��6�l�E9�<���`��b��~̝?{�/v��cbD���bS�c'���ΝCS�����{���}`��U蛄&�!�O9GaY�8�A��2�P�sk'iP�a`^�����M�VG����Y����������7{��"������ch�YX�nr���S-ZA5�j���l)I��M�F֓��4r��(Q����`�S�+�cҨ-��p��������;]��+w�["=[.Ob��J>L�����݆�A�_٦÷Y��p�5:�At"�/��5g�i�?���L�F���ы�u+�M ]�S�f�`21m7 -[ӽ^�jJi��ˇp�:.x��mn���&l�9��_�b1=N+{��?�Tq"&�9�D�"E���uxa����/n��F0<1	m�wߘt��ݙ4�5N�F�͉��6�OЖ<�k �����F�TI�d,R�4���xu{$����8��c �M�
�=mi�Bu�l�CN)�NVn*��E5K�8|N�cg$�@�����R�F;oia����c`%,7_Sc�����XG�� aŅ���io"4ߐ��+]p�I�%�
S�5/�B�=WBK����Y���A,3+���)H9��*�@:�IVހf��C�t�_�����3(T��}q�H�V��4z�
���C[��HG���H�$'<6:�M;va�@F&&Qo40w�+�+o���-M�c�r�Պ/���TG�ydӢ�Z���#���gwb���0�ߋ��^��Q�x(OTQ�zB��@3,߰Q�#�l݄؟:���[���#C{�J�nݴ�S��(�+b�V��v�܅ث
hg�yw�jf��#����g<�Gyr�C�X��k@�@��ퟍ�����A�MUR�u�4�͚���^9�!U��Qڎ8`�|�j�U�(�*�x[��P�i�������Z� ��P5�V��E2�"����^I'�4K�63R���I���"&帳q���	���#{�P�I�cj�݀��A6M�^��Qe=��R�p�E��;��A/E{�s ��� ^���#A`�RURo���W	���W)�8Һ9�x��=1�j��eK/�-
Xb���\z���@��p�*��si��?b�r�1��h����ZHs��6�5����"�F�g�6�4��8��6$:��m�}��"A
��^�m��!�%�m�snJ
&����3�ew+��� �I����)&>��-�js|7��g�%@wg�zAP�$R_^���{]LUj�(���:1]*K��do_�8i�Ho��/�D��p��Ճ�iB��5��,�
�Ue�r��T�G:�M�X%id�#W�	����VH����P��ڰ @����`�HmS������h	��@��c��M    IDATd�"�	M3ǵẶt˸E�X�\����
7Ř0��Ć
𫚋F��K4��P��C�fH�sU�����f��В���@�'Rpe�)pa`,7��j�1.�R	Fցa����	G+��~`�p��!>i/����$�D�@ã��1���(윳O������`Y.�5�M?�f4��� uˆ��7� Gs8�z����)�Y3��PP7n��yp��|��믪��-�a�┖��y�����m�.l�>$_�A������S�ܛ��%t�_��KwÂ���混d���#LԂ ^����dpT�>�r��!P�$�[QR/�ڢ۞Q��qrڳ����V��L���B�f�
E�)�z�:�4Y�=Lg;]Y/���
M�.�^w�*�9��+9�̗�p}I�0�@T2��ol���RC}����j۶t`��n|�S�oY��j,�_�p����S/n��D�����Sdo?L7���e�X*�늯o�v p�V񌤃�kW�Cl��{��J������	D���'
?�$6T��c���\��+�a�%�$��d�=���C�C��TG-�9'P���ig;	��D�����x�oo`gӑ�?�6ڴ�ЙQޅf�Æ|��b��`Jc&&�����'�T�>����[.?��<��ڳxm�Rf�t��C�bd��u�v
p���ӾIA,�a�T���;73��}��*�PH��� �dX[[��`��Z�����B=X��P�,17�d���dF�DƞM	���EKG��6��$��Ɛ���5��b�n� �����eK�O�&��ڻ��k��-EF~��O9��S�Ig��Y�"L5�;+1lM�ޘ�Sl/���J�<15%���s�z*0\��m*jhJS&aZ�H�nz>
y���	�X�}sz1U�W�%8l�>蕪D.��ɒ�Y CUR�h��~�N�bxt'�l߆��N��f����H���E�F�\��oegXP���D����f���E��	-T!s��K8�-[w
�!�A���u�JJ��SOȱG}��>}��`�\C�Z�����k�rYlߴqF��Ձ\֔�Q���D,��3m�<�^�R#���DU"�J���'�	�?Ӧ�����̴l��V���j�н���o���C�ьjS�N���Eii�i��-�B�h��LA��uBcOEz��.҅Nq�r9d�U�X
Y(elU�"�ڳ&����F&1�7�/~�~�I���+��z)�C�'�rN:�v�1x����d�5{)z�`C���N���-��U��.Z�}Z�ժ'�H���d���mӀ/�`Ǭ�FQ�2�1�6*Jny��ڱ$h�1u�[>��!�6]��{�|��K92f��7҇F��$�u���B2�+��\KО���].��z��^Q{oDr?�;�[�7c��>��+�T%��E�[R9~7;�x���FX�`w�cₓ���U�X8㈹�::����.{�i�(�a���=��T�5�6��u��Q�i��uԔ�uC�T��4+�ؼ��,&H�n���`i6�ahh�%�J�jPQ��RFȢ�������B��R�"�H\���=	��5��t�� �E�c��o`��!"m�͟]�a޼٘?oW\���=6VF��ڂ�S���ːny�\�s<�/�k!�5�J���Rp��I�ba�d�T��xm<^�R�fR�7s�8մڬZQ �A#�g�E�|���Kȼh�\��q�9yS:�m۪TD���y��+}t-�(n�ruIbg�6�I,���X
���D��S�Lk��㣛�e�vi�|ž��������J�K=6�S�_�n�y�	�u���ts���,uT���,�Q��X�'�a�Y�v�K��f��ў1p �l#ۀeɊ��9������T���}���W��Vw�pN�
���7��h��c�R.��c�E�����a�LN O��˸2�U@�M��J�"J��\��Ρ�kw����1陼���ɠ�+
�\I ����](��}|Q�#�Pc�F[$��m.�廬�D,���]���w1h�>�׼��z�R�G s���`�-�7���P�H��ΉH<�E2z�\Gv\�5Z�+�v��[����$�6��\���Ȣ������3�w�{���9�<~���{~�����>�U��V��H;���D �B1ˉ�S)mhYh����YE��"(�Ly>x���b|� ���l $�	��O#5�M������3��R��aK��`�?�?݇/~��w݁��)���Ѹ��8��(/�$���48�JŁW1b��Ty��W:X
�:1�n|�/�l�A!$�C}O��t�m^8Co�8{�Q�p>��[F0�Ew��3���>��z3-öv��d,�,̻T��ᥳK�8� &��{1�=u��+�q�y�PA`��`3��V�d��
�wY��(��]������H24�����w��� "�*>"E�Tc���i3S2���`��G[X[�㾻�ŷ��n���n��@1��K5<�����|��*H��Eg6�͉j[F̲���)�������"~��S��bptW��{�n�ܳS��^�NG�>�'�2=`1[1�`�{��}]:y�o�y~I~.��A�C��X���D��Y�Pq/]F؉!䨿�l�Ƒ����P�-!�@6O�	-ɛ�ͦ'����D���j�j}ف���Ig�=qe~I���s|��y~�LZ0�rm-�~�I�D��\7�ťu��.j�T]\l1@sC��_�,�t\62�Yq�B�F����#R���1�-y]�q���Ln*��QO����6��J����m�G�7Sԣoȵ��&ÖɆ��ۛ ����5�P��Q�w!�M�-�}��`ok�5ض���E��_z�x���x����2H򲁓����Zƽ��?�Ǿ�'��/���x-"�L�f�0Lբ�ǈH&��������+���S�o�@�e�><���\�%_�>8��PW��h����M��b�B>��%�eT[�<�l�C{5Y#��&�� �\�OU��F�ԑ2�29Z��n8� X3:��ݑ�=��aSs!I�u��Э�n���]q/g����p!���ߍ��uܷ�R�c��x� ���f�kS�(�2>�5R�_9����1E�}������
��1tM6�!�,��4�{��p�������e6%J^��V�3�$��ʂ�����]��ڇ�+�Gq�dO�5���E��طg
Ŭ�J���Nai5��tkt�1��;nW[�L��r�2��/�į�����瓠@�i�c``xC���4A�C��T^Ǒ�^�r"����(�\��Z�vj�f��=ϸ�0 �:�^?I���5"b�=�`��	�ԝ�F����4Tw#�6�p�ur��5�X���B�i l�p��nrI�$9�%E<����PG�N�9�TZb"�̜�9n�ݸ��Sh�fNu:���_�e21�~$[�l�n�G�`���b�E2���82(=r2�h{ǲ��n�^�'�Ɗ˥.�#��M7�F���׺"bU���Ҙ� AW��f�\�"
LHe�g@����>�JA&��1C����>�JE�Eh��d?���t}�O�*�E�ôc�����p?�y�f5��k����&R�0Y͊�6t��3�IԷf���c�]+i��g���oU��'?�Np���G���o�D�ǾY��=����~���*��h��Q�)Y�U�mXf ��jx-�`�#�fl��5J�&	W�yȶ��=�f���ڐ{P<?���A��((��Y���D�ؕl����a�j	++u��3��ެP�o��9?3������J�g���f���s��r�+��SՒQIP0.{�_����C�(�m3��w:!1"��L�p,8|�!�)��k�%�%�i�d��!Tx?�Z(7Z��|T��z��8w���k��,1M���2��>���o�̸��=8T�9pR��]�52��t1R�0
���lT����R+B�8����2������6dR1�S�E���ۧA������0�u12N���M�ϗ�|�L����Q��01I�P��=�u&����b"Nõ4����/���9��2���)� 2zT�7A��5�L���4U�4���Az5�&k2�b0k�Fv�e>f�r�D����
�qZ�;n�"2D:� ����LLk��'��������4�趈��ܿ�0RI��"i<�)�:ڞz��M�G�->���B�A�@�2ټT <��WK��"�����ۀ���ܵ)x�V���@�$_=�Z��W?
r�Zd�7ez�F���a��+��lҢ��5�}4<�T��Y���Z���$�"�"�A�����f�!�íE�~��Ű0#�7'�T�J4�2"�lfL�=fw�"����B��-��D���{I�.�,��]E�_�}o<�Ǿ�-�n��uv��)ǰe���-�Ù3����� ?xju��(�T\���m�D�UO9�ײp�4�qC�	�ٴ(�+D(v�%$P�6mLl���I���2q]E���h�y%��1\�ENձ�65�z-����<{'�\��S�o��:;�& ���KA�8����|$=��8�����0����� Wņ�B	8�d>X�e�j��19��[��_CE���S>sn��AxiR$iiIl��w\/���`GO�B>��J��K�)z�}��+�����`�-7�A&�75���k`�Û,��ő��掩%[�Wԉ|d#.#bs1�iY�jvɌ�C#"C�RǠ�u���n��]g��E:E��8��:%�=�m��5C�c��:~�֫T�!��<��h7��D��H/.�j
��c�M�%+_\Zę��15�I*�Aa�K2�4�a���w�ك�+K��������+�)��a��ז@F�F���(�eY���y]�gX[lIF֧�m�F�V�o�� W��#��P�H�8�M�Z]KF�,9w���kp3��rd@�I���?:1�6�1f3�0���eCfu�3l1��^L�iGF��'��#���f���k���������5�M݉'��&�0:� l���=�tġ][��P-=�A���h����S�H��fb��!�࣌_��&�ƋD�g��D4����CL��ĪW��59���| Ih�FUѤhXo���avg�
��o�H��\�D6�L��e\�g�ow��Z�C�*��%�ʿ{O=�~�3�!���s5�����T)�@F�K����������Q�UǢM�q���^0#�8�n�*V[^<�J� �#�&?��>�f�3G��+�O6��v\�"�|O6�~!�B��d"Oʊ��8-y��� \㏙I�P���dK��������L��i0��%m>�#��ro�eY������V�ƙ.oZ�N*�R�)���5�05����ލ��D���(��A2t�m��-����ؾ}t�HM��q6�ߗ.����<�D ���`q��Q�a��F�ƖF�^|@v;��x���TS���ř�9UH3�����e�@"��é�%��%��>�X��J�N:��֛�k���L����ϰ<�Y���K��Xɠ��~'*�:��p�}�C����^��/i`_X��qSXXi���ٹ\Y�Ay��$�P��dZ<%qq�*���af�f!\�>�LV�:���"e��Z��Ds��'TX#e2�}g�������m	i%������:���v�e�^�b�T'�~`#n��GG�U3���r����$�]�r�%��V-���oC��÷�O�\[f���x����z�"U�9ˊF���gŁ"�#q�!m޲���>�^�J 7I� O��>�u��j������͊�cZ?�(�H��ܰ�������0�k��M�.�ۚ�Ȯ��!�a����y�f��z��= Y=�-ĝ�����ɱE M��6x2jҠ�����J�H����m����>G$�����n44�>�F��g�m#��ѪwP�`~�*��?�����"��������|��h:����	�?��ￌ�oۍ���'г]���d��V0,T��dV��p]~(����0B��M`�f�.�iJ^0���9iK��/�M���?�����_�w�4C���S�Mp�6z��u��XVPC�	@�b6�V��r=��Ϝ�*H�2bRv�� ����e���N �$P�^w*�����B�S��X��5�%�ۿ���;�t�fs~�����:�ˋ�KX\\��=4�Ĉm�*Ӏ��5?�A���-��e����	�/�|	�~�u��������(�YȲ��$����>u���� t��&�&�T�8ho2�L ��a��(n:8��Ɍ��m�b�" ��`��y���Q؁=,��c|���%�~��+��s'P*5��s`p/�9���~��H�eQk��_@�ۑ _m�6�C\��&\d�Y�����1]�Ӝ�ͧ�W@U3�3����س�
ݟ�����x��{C�	y��c����X��%hs���$`�H �,�NG��R�Xb�C��t���F��5���U���!���B�VCz�3h�Y	�Ն'���ղ�(�ɇ��H������cS��T�
�I�T�왳�e�.��"��D�;��K�q��)���7#�) ��Ȍ$��y8�C�T]�^�^�D;���HA�A� �T	P[%����x]6u=��x�ik~�_�����PQ���z��}���&�%B$�l�Ҫ�����9�A_;ܓ���)��[�$��YI34�P�Q����h7�ǻ��O>�;�J��@�H؆�C�����	�էq�wab��/��/~廘ڵ�K�`�;��%���ΫxvcH��M�JC~��'�Җ��"�+0�b�ѣ�U����,���Z�Q�[�t!��g���	�4b��n�M�?Ѯ��{���3DJ@�� ���3`w��xT+伮o��O�'ʅ\D݄��67ˑ��u�ß��L��DS,uQ����N1k�=�o:�� �T�n���@k��<�Ԩ�pq^���л18�V^g��b��ݾ��8s�fϟ��[oEz�z$\��<w���\́�Ž�Z�,*}f�����A"+B�b��/e���RR}�� ��Ǉ�S�-*e��e���w߆��b2�L��N��w+�zdv��|̟[AieK��K%<���0R���8�f�15=%A�՗Obe-�а��/]]S�Tި�1�N�ǟ�ha��dK���~�)��O������[B0�I�4ef`�o�Ϭ8��z�%>�,��6���m�6m�+�?7:<�d2-�Ak�k2�fG*E��;����q�:N�;��-�1:�p=�x��a�!	6-4�D��&5I ��[}t;��-cf�$^=�
������W���\F��0C[	�+,^Fye6i���c�u���T(!���������d�pc2�|���1w����Lc�M7I���	$���"���m��	n�T�٪��7��cmH?����#+�����Q��`�-	�&��}-�*�4h�2�hCy�Hkbƾ5��|<���3Xsq>"�M.8��4kf:)[�y?	��Ez��.( f��m[�����:�vl������XY]U�����������ˣ��'ލ�?�$�^�">�	Mn4'��"�`n}�au=�,����RQ���g����(����&(@�߆%\	���;��)���j%G�/	}�SE9�>�X(��~�`�S`��4�`�J���jC͟�"��N$X��2޿���1�N�ˁ<�fn�$h�R!RI����Cj�==jԒ�[C���@����^�����n����-��$��ȑ�044��s�f����d0��3�b�Ν���E|�_��/3�'�ۅN7�@6��}�,��G�KZ�f���w�'�!�>�)-�,��GG�)�����RJ7����F�]t�E<����~�w>t��\���i�q|��<l�x�W�����;z
��e�;n;t�V��p+�\X@:����*�G&p��[�jy�vX�_���!�p���    IDATq�t�5}Y�d�=��N�K|kZ��� )��1�r�HGt��<�N�5SׇX����ʆ��ӟ��A�#�#+���������Q�~�V���-r�j�����_r=$ �Ĭ��k ��1w�N�>�~���=7��;���![@6�C��A��1��<�n���e���@Ŕ�{�m�vё �sn��z�-}y�Σ��X���O=�T.�ɭ�X\)ᮻ����FFǱ�^��jEZ6���C��fuO?�)լ����Ʈ]3غg�8�Y��4}Þ|�9k3Y���Z�}��A7���$r��z���9��4�ѳ�����0���L��i>f���O��4Ѧ���V!�EǠ0�/�Ǒ�&%Xи��������	6\b��&RdVI���E�N��zM+�~�����;�/�ض'��s*_pu��Ԥ�����u���� �xOZi�� �EEEI�3j~�BmS)��)�?漃-�f�.��|6��'ID̘s��$�T�(S�1	��R�^>>�:�^�h_k��ⵤ�4]��N ʅ1߂�p`W	��oxD���1(�ftl�8�ġ�����/��:���ġ�
!�zݏ}!t�\��B&�i�α�� �W[����0x�-�!�]E���o0�蛓�C���O�^kahx�\�
u"�8s���:���������	l�>��4�_\l��p��
��b�ߨdy�$2�QQꓛ��2�bL*1��L/.��8(c�Ȋ�rR�qZ��)ك�N�E��&�Ɠ�������{&%�nKv��H�A�W�2��'�|�;��±sW�=�<j� ;�'��|l��F~`��z+�ƆQ��00Q���s����+Z�̞+� R�@)��$ԏk��h ��ǅK̳�;VG^W���a�+D0��M)�kD<H�K�ے6E�c�լ��:??/s~��͇��vq��!�����[2�}��*3��T��;�������19��K�ӊ�-&Qn�BX&3Rrl+�\��}
��Y����C��9�� �M��4�.�[�V��QYC}eI|+/^�"?�\##C8x�ر�z,����l��	ߓ����%,.�I��Ҭ
�;4'�x��ߊb1/PC.����Z%��Z_�Z79x�L[����t��W^��{mT|&ێ���_��)��_.�3L�5�S8�1[�)y��=�kN�:`���dF��$4f��&5Z&�����Y9����F��@^@B��z��+��Ɵ��O!W�D,ђ�}�]wH��g?�x����w�Ó�稯� =�A<c���JbR��o��MVc��ղ�.�ұ�s&S�I�/�W��03#�U6�k�
k5��#a��1'>�-��I?�����O�����X��<[̺�xN�O��]�y��7����]��D��~ρ+$1��l 1~@�*I7�u����:��$�J�7I�o��Կ��_�W��3�~��j�WTj_|�TǙ�	ڥ�j��P��ݏz�l��®��p��%x�����r��d1:�f��Ϟ�K����x2��C�O"����4�1}ѱ��jfC,ii(�5r�v�̆�8;$[0�%,���K�pp�n�i��E�l�6}z�)����-y��E|�oÅ�� �v_�δגn ���Q�~�F~�҅����q����-�P$�V&X�  �QYԆZ��﹂*�1�$�NB)��������-?�X;@���X63����U���d�A�t�.v�݃�����"�
M���|L��<���<o�Js�_�䄶����Tpˍc��PWk���&N�R��8s�U�c／7�����܍|.���2��t�K1u[X�p+�e\�r^Z6��]/��u�nܰ�f/�J�!}�^<w�t�.̢Q-aj���y�޵��#r�Ya3H��ϵ^�^ƥ�T�\��6�_vԓ��[�AG[~�d��O^�K}*��σ6=-e�������1ꖮTz�,��#�L�0D�h��]���-��s�ß�@��C���R��\��^�n�^Z[�F=V�>�֯��X�o������$��@c�K+�.�����*Zı��v�F-�C'����-�R8��]�S��vhb��V]Y�w�3��}���o�]^�u��Q�=/p����H��Т���)y��4ܼ�+�lI��q`s�CMHK�9 �z6{X�mD����ݖ燶�L���W d+�� QJ*	�z�{��fr�&r��Z�|¹l4���Z%<���x���13=�L�'TdB��l�� ������^��c���kv~	?|��8]��"U=��{�o��Xa�[Ʊ^�^i�6�~�	�Z!�0��e;���&*&3�P�i*������f`E�^|�F(�p�^�}Jfw]� ���=�ئ��	7�8�D��z��(�R�4�a ��ǟ�ٳ���˧PizhwzR�p�i��zLm�"���n�ԋ��[��f�&C���p��c�.j�*0ñ�_�r����,�ڮ`���E���B��m�j~F*5���8�Y�����g�����M%QZ[��'D�AV��i��M��X,"��J��ߧ!A���(b_�_�����m���abt�mن�������XꅉX���R���������u�<�毇n�Y*	�,�W*r��8ծ��8���%t�>J����Ø������@iлV*��^A.�F>���?{N�S�jl�#C(�}��yOrX���F���jk��X���Q�c�v�
�0CG=���
|�f�z������W%6��0�nm�h~.-2)�Ⱦԍ�����Yr�:1 4[Mٸ��8����e�ENVX�y��B<&627"IM ����o�ICtaGC�ε���c�"@�ZǾ��x�����d5<��E���H�.ݰx:�:ؾ�V9�����L$-��/PP��T� yn��R�Y�v��Y���c�H�x�붣T�㙣+x��

9f�>�������>�����Ou8���N�(U*�%���6ޯ$�p�
�Er�R}���$..��C�M�}X�W��"'�b	eQ۬OwVN6;dJ�h�v�r))'�F�G��_wZl�N�O~��pi��}�
S��E��)���3� �=D~�ʅY�,�pa~�/^��J	�CC�'�B��D��� ~���߶U��-����3�[(���:z�9����G(�N�'��fD�Qe�JlE3�H�����5Ўܸ-��
L��}��p�=7�Pd�TC��3���\����DXi����<��Y�LGl%�f�ؽ}�����(�Im��c�1p�un���*N_@��:M���&��|d��~�j�%��l�U��Y23sҫu����lf:ɏ������t}Tje�c��r�?s��V��������8�N[�l��SiZA���JY�f�4`��G�\���%��s�m�f5��ST#�I1�JS�6d���)EYE����˸��[�{,��'&��f� dK{�:�ʶ<ΚTW�a�������&�5A`�<���5�R��Kb߾QSYV��Ɇ��7�� Ui�K�_����wŢ�����&�?e���
�� N\UDc%'��X�׶O�붑Ŋ�[�8��Cd�mo����i�Pdhh�7�E�XHKdE��+s�8?{	w�vҙ��8�DiA�y�4s��`�3
ؑ`�~8]B>�T�#+I�ޙT�k[h��h���oۃ_����k?��E���|���,pٷ=�&���=�|AW�[�ޅv{	�v߂zM�l>'r�\�nv�A��VsKK�����u�����}7����o|��Ϗ~�~�����'���h���-(�	�H+$��.vYb�V�c�O���ėy	#|:�D�ۅ��Z<�cfL!!����2���<��c�����K�`{��ڞ��[o����w�>2�$jkm`��ls,!�ia�u�������|�������;H}�F�Ξ��+�K(/���ŋ8c�/�/���!�J!f�����7�û+<W����f_3?x��}�"*M� -'/����.�'�V�̌��7j����'�@��ۈ
���%�oC�۽���_�ް�LB^�*�fIJV@�Jڛ���o}�k�_,�����̒P���ۮá����F��}���W�	�J��ᬔ��K���v
�׌yh�ݧ�=�DR|�𔧏���]��G+� -{���o�u�4u�aiL$�(b�e����+8s�,hPq��C2�ɐїn4:�כ�"�@���� (� |�4�E,\9�Ç@/i!���4�P^����.�S���س{�VEc��b"�D2��"�4���3Y_3��P]8����K��&&%�K��dy]q[&�}E� �ɨ+"ρC��sr�UX(�p6 q$Ou:t�Q�t��^�o5
x� "(^t=��-�����	����Οc?���l�Q��zI��=%�h �}-�lÕUB	+!f��R���Pl۾��'���>n�� �Ǉ��I��Kf����е#-m��=A��:���Of��V	�D�>�a�A��zYc��Ç>���A,����wP���������~'����~U��:���]w���5�R���B&�a�n �T��*W��^�f��{p�M����9|�][�2՝m%Q��08l�v$�Z��o����y���d<���Ռ3�⨰k;چK��3E�D�@ZZ|�m�,[8]J�	:�V�%Z�\��h?�A"��K�ĭ�>���F�-ψY�t�=	dE��bυ����5�-��?|7�r�A���O��N�.0	ڄs55}�[ߑ?��W���WN�ʃ�]<�����:-�~��PH�n�T��p9���_Ri׋�M�����8K�H�4 ����T�XZeCgI(����&�K[� �%:�0���{/��~[�ds$Sh/��>5'ԍ&W�p��%���9{	sW5{;qqNq� ��*���;nŭ�����2F'F�!�ǯc`�:�je|���cb��h6��u��tW\�g�;ys
���B�+�ϔ�i0+5��P��*x]��o�kDO���eKP�v|)5ɨ˲�)�}gC͑�ꁼ���Ed�)���Rޕ�+Z�Tˋ���m�z3�kVW12�EZOH��Iw,�ZW�Od��2$�=j�d��qG����[Ƒ��ɲ���h�s��k*�R?�B����ʭ7[�W�}�`L��@<������L��-b��d���RnV�w:�0�(y����$2=��StH O~NP@Fg2g���5���o��PdbȊ�ص>�P��%���Q��Z��̚��[�/NV�����H�m�_��G�؉�������Ɛ�	a���#�q���L3����f�O(���hժ�L��;��ؾC]����<��x�#o��~��(�T�������'�k��s��w^�sϽ��;nD�HS�k/�f!��"K�F����~�ޏWO��c�ݎ�j]����Q����/`���P(N�\^4ɗ���J�����ڲ��i���2�Aߗ�ML7��|>�!��lݬ�i=G�#�h��nZ6k��� �Y�,� ��'L8D�F���>3�lC����{�ny���D�!`7���(���0f5Z�H�C�w�~��>���pq�Ǎa���A��f���˗qynO?��|�x���VQ7ʙ��xq�#����n
7�ۅ7��v�<�%Y"��2������E��XM
�^����W[�)��*�T�F���(�=���@=�l���S3a�~ő��=�G�<��2'�5��;��ʦ�su�������~���9v(��]��'q����;Dg��{�j�9�r�tT�8{v�LL_�z��C��\�6�Eݠ�Z��\�vn�8����5Ȇ��mмE7B$�����FЖ�3&sS>�u�:a{�}^.f	k�����݋��&BR��D��{���$䐋��\17Ϣ, 7�$��
��'vc�����Z�
��n�l� ���ƅ>��EM�j�-�|mj�����,$�XK*"ʫ��Xh2+^I��(�0�Þ�/-F���
c��f��+�$����8q L�9G�Ԣ�E�˶�����u��'�?�T>9����Z��Z;K����g�\���"Ny¾rB�"��a�E�j���9��2�/q�Q�C�y�=�"�4e���.��dd"��P�M�΍�:�zd�)�	���ȉ�B䉱�+88O�P��5�D�A�ȧ�8|ߘ�!�Μ������
:�s0d}��t6�/}�o1{����t;~�d��,�mm�~�>���ï��~���CX��������^Z����R�,��Q[�tf��cx˃�_��{��\A�";�Cm����S�1�C<�l[D�i�mTM�Ie(���Ik�a�g���y�*����� w�+UQ2I���=i�qY�{��e�O����u��a�F]��T�}��nS#�]S�J�FEw�Ņ\�� ��_|�O���Z	�6��օ�?4:��215����^��4�܉�_C�L�Z/�zA��+=X�� Q����؉�>��ADF�Gyr)�*���v�/hN�Y���/>�����A��5�����F��cmL��܂�V(������s(��X\�>o�V��O��O���˸��;�m�q�Y+�0{�U��.aeQ����2J%3�d���w��s@�Ǚ�133�s/�8���K�a���a���@)�Ϣ,N��s�F�v�p>C�5�H@K�M9g�"W@Wn�&h���X.y�z��-��)$A\gB���Bl2!��;�C��x���11�`6"ҹ��M�%*ީ�P�ĕ�B�aZ�0�8�e�K�-%i��:�w��?o)U5��D��abe�@h����Bs%h3�d+-���&���:�Β9H��)rR��ֲ��f_��H�~��m�x�5t�
��mm��\�5��!��<�F���e�Z��ٗ*F�8�T�:�����W��ז���sr�n��`T2c��^�9VM<&f���z�ᙠ)�JE)���=ԙ�Ko[_gma�F����-�*��/af��];����O�C�<�zT�������ϩ6I��"N��؀nά�b=���C�� ���Զ
�&��".^���K�֔�/�w�]����"��o
t�;}�
�?�'_2�}�z]Z������m�n>+̪c}��MX�8z��Tr�x�4L���u
r��	hW��e�$�sҙ�m.�N�a,��;IR����WB�q����4D�!��|���a��i|��~T�N%��l����ҥY\8w^n��g/���q��,.-h�y��2��c�@NNMb�P*µ	����D�XY�(=<���^^��:q��_&��-�(K�~G�D´W�N���fh!FV��d>�A Q�W;(�$�t�t�ŁC;�c�2~S�K����w�[�)UkXYZ��bI�赦>��KW��d��)�޹�Ú=�q��s����'e t�c�����1l�mI��-�t����ѩ�6�)�����<�8���Vjfz�$ߌ�e��ju���4e_���3(y�P|@#�%}H\�tڲ��	[Ӡ �YZUO�
�}��/&��M�z��\B�H"`?֠��ɞ:m�U�4r]"}Gf\�;<&B"�@g�#���2���6-
2��J����cl�$Xۮ��z%Im�!d����H%@�1�&����P���i��0:�S�����A��MR�%FP�4�^�v��B2���\>}n���(�PH'���O��� �XƧ�E[!.�^�Ν3Z���!���tn��10�1��-韇Hų�]vD7�8�.,�`z��2P�x�m�P�	�j׫��m�05YD�������!�\��'����;9�����?����<�?�ï���
V�,A��A���N@�@������#c�4��s�ȹak�13��!��L:�L��࠺0p�9���WD�_�c�IsO�m!�Ɍ�{��>��i�����|�#Cv���l�.�S��%)#�%�يn� @�B�[G,����Uj�Pc6a���p��X9����l,n    IDATº��ڎ�R����Yh5+h�xsWp����_�(�}p�1�n�ewX[^��c'0����g΋����k%\���d&'�Xtg߹{7n��&8�>XC�,��$����8�A�85�㧗��K�t�l�8�?�t��d�ϖ�D���V�޺&�IF��i�]�62CqP3�T��<7R\�P��s��1:V@ק�E�r]2_��RU��W+X_������?�1��o��LR��^ģ_yT���Tˋ)�l}�;^D:��d�g��	��\���`w133�d$���i��������X���`�>8�b&o&�-�#YJ��j����X:GP/`��LL]ɨdfO)o06�[����#t�4E�!NH��@��vԛO��T�[�:�`Bz_�\+�
n�����:�x|��|�)1�r��%Y�q:h�	����ض8]��S���sn<l��Cy_s��8�N��M�9��M?�6Mhu�#
�T�c�b��}!�;�4��+r�7�'�dZ�]Q���I��%!E�����9R������N����.f�BV����&<GZ)��"KR)���j!7J�Sf`t��B&�V�S���0��3��[��l��k��p����u*K�ē��>�.�|u��7籼���wLcx��x����>����}�v�4e��bjT[[F����~��������8y�i�X�qL�V�Ϝ��QkjBI0¶m��g�.�/�	}����#褆`%��2vjT�T�t����9�=E��3��X��A�SA�a5��22PE�n���	��X1��by�"W�\�w�Hѱ����Õ�lS*f�)���1x� 媪���)����059��!��;������8q�$*�:��k�zu��	y�x�Ɵ��-������Bqz^�f���LI�}츾/w��F��U�_�>Gr�!opz��Ϧ`�	����`d�-�D�>����1���R����p������b���]�q�Af%��R�������s��E��F'�b��U4*5��;p=n��.�W���Oj � ��_�s\���^?���b� j5����d�#B��_>�(7�Ze#C䋺i�sH�2h3�"��q�-���XV�#��hhF��f�3m��j�J��( �5��l����7qv'��g;�[��w>-�x�6�G��k����ѠT�4�H)-��)+9�bV�!��<�Ё�f4~O�g��&�u�m�u�W"C�N�Ul��������χ��r���T&옇����%+nj�3c����hr�����{�u���Q�H����F������I1�̺��<�1t�&��DAON����ZDD!GqnC�G�UE���C�{j��8<�#����<u��� tVq�Oj$�,�$�M&z��jǴp�Ra�ƶ�5��r�*>�����<�ݿ�?/�����(Vf�HRh��驭��:XY�8���{��`!+��UxU���o����A��G�u��חPm��)��(�V���3�ᤴV^���"��.��=�=3������/���%2豺���DK�h�Oz^�-�j�=:�2�2-|�#���G;�ʱKػ[5m�|�^��?E�~���+�C6�B'?.�"ü�������=��0�#.l� ��Fw��F�3�SطZǧ���K7ܰC%79�Ivq挪��8q
��]@��!�Yx�E�%-W���Je�����y�Nt�M��%$����b�̌4�[f��ꫳطo�=�*Z��ݽ���T$^?���[@*���.�w1�f/S�K;#�I_�E�l^?]yg��b����d�&�D��QLl��/�V%����jH�X]YC�^G�Ґ�a��I��G> �s�Ѝ�ƻ:�H��S���*����Z���aHQ�q�6,\^��%�y�7�eDZ| ���`�;{��A[jB5J6�-�W	n�~��;��ԍ`6���Ag���J����@�:����2�#zG7:�)��QE�DƲ�UH��и<��*
%��j����C�LR��zm)B�:+��G�hFco�.FB!��H�7��P�����V`����t�q��&�U��Pvꨭ�u.�e"k5�pɚ�!c_�XT/[�|�E�Z�k�?3cX�xfd��kA�>�I�wD-�ma1�]Jߟ���q4��&�F���%uy\gi"�51w:���<�{+4�ةC���~?;���
�k�Q.-������o��޼���?�����c�{/=�����;�����9�?غk�zEZ�l_I���O��N}��9��W�ǿ�qq��_:�v�.�]Q�}nX4�&�S�\]D�19��tQ2�g��ş��7P��a�t��dZ�a�ѝ�ή�v�^�
t���^�ǝ������{�
��C�$�z��3x�x�����Q�Xf/.��u�B�D��vj���$��76w7��ka���K������'1�.Ȓ�,�5���L����� �r��{�}�4/V\\?|���:�"̥�e�_]D*Y���� �CC�y�N�k�2���o�-=���:N������va;.zH�o�7�
�����X�:"DI3C����f�B<-��W��'5�9�%-�פ-��~�B�G>�A=�E�6���X��Q���瀈����E�Qk%A���Y��0��ߏ��i\7���zs�.�.�� ��c7�2B ���hO�RV��fY7�t*�vXG<�B����`2����"
漃�g��9Z93-�,�2̸8���ŕ�dD�Oz��;�!�1�k31�E?R\3����fغ����y�/r g��
md���Q%���av��a���g)�~��Dcwm���ϦY���8X%�]���>0u2e����2%E;�T3W1Df��+���̇C�HT�HWH9�7S�}�><��֥��,R�CqB��(��#mT^S1���R�%�h��~�a�X�j�m�vT�qs�f��zn�<N#����d�g%%�5�+p6H���#x)�X:S�r��j�Mضjm!K�Zڶ��G�Ǯc�����9V��߾��������;�:!��rA<�B6���:�W�ˠ=0b�֛���o܇��4��vwU��D�ڷ��������r��輮Z�bϮC$�o�����^E'V���
Ϟ.2��0hs."	y*��ܿ17�>��_�'��ػ�a���q�����$[������^Y�sϟ�������y���m�vۨ��(�����6۳��G�R�5VO^0�\�ϲΑ�B����%Xv{v���;��#��F}����X\�(4�;�ť8y�	�G�_�gJ�-���ɏP-�٬�czB��cC�8��Y�����|�YY�Z3�0�aT&ʍ�R4��w��q�����]N
�*ur��4N�]Llj/���5Z���H͎�l���l��.�Nu"J�.f���#�'�axxTt,�h�{��}x���/,\���k8z|���:�t.�j�����ɮ� �@�h��h ct��e����Q��(��m��Rп>P�s`�O)�9�A� !�\�b6=dr��$RQ2��:�#����Tʍ�V��F
�߻���Qd�Ș�����#S=M3O��"B��!��F�_��Y���S$��(�jT4�(-w�}��:���3Z��N�A�m����lA�+�Z�"�e$��B!�F���/}~~'H�2XgZb�!�� ��#�L��G�X|��J\K��J��*tN�I��l���c�?���3����\�TBr�"M�us��FZt��Scw�k��N�ehZ�24��j{�'��Y��bb�\Z+��*�k�h�8�n#�P�Աo�V|�#?��:m�yz�G�(��hUR��w�F<e�����
^~�"l'���\4�"��ߴ5�����|mˌ���U4[5$)�A�g$�ö�'I�N�Ɗ�FGGFEi�u'N����5T]m�Nv.��㽮�3�'ZW{�dǭ�t����	;v��~R��q�q�3��2i�$p�s$��9D��,�}Z�9�pA�ӳ��h,\��B����k#�������}�82��t۰-�2e�!�Lf����?��?U�H���W���}��e)�Y&%�Y	���)R3���@&�\��,/���%��Hs��E�bDE ��ɞm)f��1�m4�%�F϶���%Ԧ]��ќ��7�E�e	�vK��`�$њ��bd�I.~VN�i��Wh��|��u�rH��w�^�J�x��@:�૏>.�UkpZO�SR���c02�M�w'.&f<��֋�b�����<l��i[D��p.��� �9����(g~� 4Dw�d��91�y�-"�j5����N%�V��L�M�Κ�iO��qɜ��7�B�Ț�R�Ak��`�n)�ࢯG�H� J+&�(�.�s�mm�?�m����3콛>tT9�-�F�!���fྦ;M�N2�UVW���@��H�1�N�~�q�]�gC,�ѿ&�H���!�p'���|F�)�]����￁��*R>y=�ENm�:O|�2�!�٪�4�g��I��!��s�*��l�F ��_�ܹ��b�="��1kcu�
��,?�7��y�e��/}Cm��G?����G�}�6���p��8�V|�?}kkm�y8$�H"������Qw޹�|���|�[�D�׃k�p3�az�,Ǔ֑'L�m�@������o�מ?��^a
HdDV�L�l.+dB�����U��`�Lo:|;���it|`e0�Kr�3��=��-0[7���H���x��&}���|=��t]�+�ny�a�r��h�È&��-P�C�VU���$��6��R��}7h漶^��Z}I/���^TQ�&��,jr-䧆E{�C����� ��+���/���L�i�>�dQ�zܮr��$'��(hsp�H�M6#%S� o$f94���}S��ڎ��l��Y=9��;��X	�#�B����G�HS]Z��\�����M��<��f��9�͞ϥp��2���#ًh�2�!,2�XB���3�d�э!�b���/�n<�;(sĊ44z��2��@ioК�E.����.A?��V�xeY*�V���<�z	��	��i-�=�W��n���t�e&Dx�4")<fÊ���,�#s����Z�G^�1�=m	1��`�"E*����TDL(���h�g�)+ AT�I��+I�O�2+��c��̚�@ �\"n�6
z��� �F��'�vc��64��8pe�4�!q &���XM�}c�x���-�B��ip�$|�l^_���7SJ(��m�u�}"� 5pt�V�c� �^c�I��d2��2��,�̞���f�o�E=�ߺO��3�������l�������G����N���B:SP�;��O.@��e�*��������νY�9e-��CȐlM����p����>ߣ�#p���g�{G����F@�^jv"%����R�Q��]A������?%��o�ޑ�����bDèM�?/� ��q����d�vX�+G+XYi➻���ߝ��^}�e¡y����i;��t�*1%��f
��ݚmj�!���I����a��!��a����=���q�R��n.��rl䇆��ZFfp3[�������NW�2�o::����ǇI��zc�a���x��� GOK.�K��n��'b��2�d�6�Wjg�P6N�n��g!��#6��V��g���e?��]F�]Be����T=�T&�B�xP�mLM(���\m��ڨ�}T&�<&��dd*Ɠ����D8��c�!��	&�Xؗ"y��j�>7]o��mɍ,Y��s`fqh6��K���ހ��F09-�y>� ks�_��^lH��8=��%�ޤ�Oۦ�A6�x��l���/�P�5D�"T�~tsb�L��8��*:qŘ�6�Z�7a��>����.?�l���R
�9��.v^�ڄ���BG朞� m�]�̶���T�͗-�F[�B6��d���
l�fW�>�v9$�4;`���Q��
X4�0�}�ވ.�P	��kĠ��Zbc63�ܹ�Q��3&9�� �~���j#�ߋ��j�ߍ#��sOR^:ma��a;�<�GF�w~�I4�x�a�A�9�P�{'�6<�]���3�������mahgR��q���B�uFT,!�dE���uox�!����櫞�5z�,���iEv����'��p�|�b���ދ��Z@m,2�Gi�df@�^;�͙P�YB?Hr���4��P2�qI}��y<��E\i����w���R%�7,�A�$'ކ�4VAv�D��l�^����0j�Uq�a��nn�T�޳����yˍcx�%LNa���R�BWW�
�b ��1�	$PGC�PDO�};�<q�}Z'q @56��]�'!2sc�&�L}���#�_���RL���'�	�\�\��v�MҨ�!p��V�I6�#��XM^tA�ݨ4��_�x��v�a����"�x�Q���J*���#&�4	eC�a�����^�95�6C9#�#Y!�3{���*���kJiCA���ѓЇ�,����L�>��ěHӃw=��,���n�9&��m��Z6]�Ŋ�&�EB����P���Q4Հ�#����4x�uX}���E�K�z����Q����kA{�*3���Y,)�r.�
	wd�C�Q���&XtnNM9�Ba���l/p)�����V�s�h�D�Skh[��?Jagf�� �{r]��Ѡ����c3�毿v���@��U]�7�T����4���|�}Op�:\�Z[<.�fX��>Q�`��G�6j+���^\����'p˭��w��.|���foz���O����Y\]\E��3������
���	@>��o��hC��^��DRü'�����"��"�-1������/�⊶�=�a�Ҩ�Y�S�ڦ�)���������nÈ�&�s�������e���_�����N([RZ7Ŵ!��DW���������p�T�x.IK����!�i���BvY
�bٷ;�>Rf��=��X��+���FZ)�,_��=�|Em�mICOLJ��[�Ț �8
DD��^�_g�I	/��("H1$EH�s����Y4d���V�=EҎ)�cT����q�	���0ڑ�L��-A[�,2��a/��!��`�%;��aK�NS���'�:��)�V�I�}�<�@<�C?G��NU,��OSP�VBe�ל��)[�TJ�a$C�x����a7Y*�asچ�O-d�t�� y��W+�n���0�$�J`S�f{�=�(j�pM5P0<w��U6�kV�iEQ�<�7���a�`2Pi7�ւi�ț���"�+Ky>�� �a��_�P��瓙&ω�v�L	#�`��׭oU	"�$�dR�m!�����l�=
2�:k�K��(��N��SY�����,�XR��(�X�y�s#Rϼh��=��2�����c�B4;H:q4��E�H�g�E���h����f�ϓV3�[on�YU	��ߙ�|kNR��Rd� 	��d
���DDEE��nD�VPQDZB����$d�+I���|��v������ObU�{�ox���w��[�4��G�0M��д��u`��'��KS\ �vBh�}xOV��B67�+_�"����p�)L�V��X����o���~�<�����/�y�^v���y�R���4�Iu�}#�-��!��4�|��x�5�Y� �=�Z�������J�i,��xǞ��`�����X���.ϡ:����\����0hl�k��v/��,������5p��o��u���g�y���cmuM��$q�ũj��q�)���s&��@�ؤ�����e|��B�h�L~љ��n�}v$V�P�t
�ip�A�M������=�3S*��hF����2��:�\�R���)�9$n<�^�`������ҩ�9����`��Ec�f��Tt���$)U�vS�2�Z�%>/�;+�y'^DK.6���������)��1Um�A'E�����=�&�r�q_�^��V���T����4�2�    IDAT]hx#���
�b�=d~�evx\��'MNX<�5\x�@��9)�{d"%����0Ӱ��$�daf��	D�~����`l	N1�뗶�O
^)���4��'�M��{�G���;*�)��;;�,����lW�EC)�YAG���/��`<�w�@��O��p���q�ʿ��E1���� �c�3�p��'EQf������H[`���[���K�[x���i��ǟQ�>mb�4��<������跇j�g��Ƽ�nx���ٲk����7[�@l��-(�1-d��y	Z�[�\�� �����o6!uG��Z���Sرc{�,���~�������o��Ux�+���h$=��ܬ֤�[����g(�vb�����N5؍���څ��=��6��t)���B|�+��K��i{�$��pu��O�g���޿�SN�����`����j���6L���XW4kl��2���D)|u����/Ź��\H�`�@)v��RXz�8z����Hʜ�[ն�����97[Yĉ��+���g�0wժ ���?��jU<֘�5vJ��u�r)+"}Lk_Nvj�+�A����I_b~�/���@���ãY�j����Fuk�v�C��!�J6_R�
�����M��aA�6��7�hR�X1%��궪�>�	�8�:�w��2���E�V��Y��BM��=�hYXbS��,�z,@m����B,�m����t�P���Q���Z�&��8�Y <�Yv>��s ��m�ѽHqq�����T��9���Xlf���gA�Tg�,�$nR3��I�����;�3/km'\��<h�����r�#�)�?��h��Y�P	��$Ț��d!t|���be8�Zp�Z�#;���7;;���Լ��{���"��L����a�dU�`�C�h007����-3։Ł��gb��1i���ڝ��|Q�����"������u8�Ȉ�$�(d(�ݿO�C�#2��z%8������A�3��K�-�VIV��d��� �1�b3��蘁���S'����L���ʫ�[o�����o��~��q_������}��Z`�B����8����}��5�P����)�wZ}D����G�P��O��?����8��}8��Sp�m����5������Nǭ�<�}�𓻏 ]2v[7c���(U4>6�p�e����6c��x�KNq� �uG6v�'Yz�V�W0���g~j��~ό�9n�@v�]�\؉��9��\0!����A3�9�TE+c�Rm�~z=u1Nѽ"������9h����,���삸��A�>���k*Ѝ��(t�.���}7sd��)��%��8u��.F��� �M�On�Y�����fTd#Q�&�9�U�e� �1��&+ϙl����T�QA�S�i��D�v��pGb��`a�ݡ�h�暪����R�3�5�ꚲ�G��TG[.�F���`����33�fh��l�I���9��)�O�Z'۞��0,Բh��^&�$��O{�}���Iv�z��	��W$�?X�� !�]0��{��q@��M��q�fM�(a���B8O�yx���t�yZܙ68a�e�A1��d�/6>��8�����٨s[۹���H�#r�I���r0�K�^����ܪ8���&���k�IQᲀwRCR�����ics݂�T���O��P��2P�h�Wo0���:�O?��}s�l随e_:`�NȨ����C�:f��0��U_���QT׏������Y�y�|��,s7���$h�C�_����sZ���ڏ������v����*�3F��5hhk�;��x
��Kaj��#G7��_���o#����������m��e�רBI}�9��F���eh7��60hX㍟'�We�Q&8`���ޥ߳i�G��2A�n6�C�e�� �����S9�ч��;�R>������K����D�麑2\����m:�E�����������7�o��R���6���ʳ9f�U�,S`՜�5]����йR��m�^�(�K�BA9��{���g����9gݒ<�&��#�1�i����s:ꨌȚI)����2���E�9ۂJoB]�lc�@��|�V�\��V��ܦ� �GM�"��YmV�%��f��Gk��BE�]��nO3{HU�3Ԉ��|j!?h�z���E!�:t����i]�"n��{���*5C�`�)�~�`/͊t����ކd<����:6�`:�i�e����(w\|m�S����#d��E[e��G�6vʸy��w�,;����}6a�P�0�<e�[m�^ȥE���x���G�!Ӷ�C���JS)q�>�r�6�l�>�qL!0�T�c��Zmk++8z��g�l9p�y(M�iP�kcsSP�7�|Ȭ�'u�ner���
�wW�D����m�
�~W������d4,bm��~{���i��U���y��\�����oy=�����~?��~�K�o�e��������Gn�i�K*ܭ۷��Xc��-�W)T��|��j$r�c��%zr�~�|a��p7��&�e�ߩ>R��SF)7�hֵ�5�
���3�s��g�7,:�c�������X>��b��.ɹ�E4��#�)�ܥ�Ue�5}���zfK3��b�����e���5��u��Y{K��P�o�n�%~�('�2�o���!Y`�u�Q�J*���j��)R[�<#%dҘ�6�.'�pe*��c����;Cc�o\� bA����DGX&�+p�J��H��@c��2m���A .ϳ��R���ck�����Bdhe���$Ϥ(kw��#Td���lL界&!ag����hvz�*�hz�τ�f�A���>�#�u �-����]S�Y;�9�<�d�PA��f�6��&���eQ6�������M6�L22���Y���c,���k'?3B�(3����$�d�!X��u�~�����.gʀm	y届�d�$a��������=Hk�CI
�T,cq.t���A��"A�)�!�-M:\����}���th��X���m�銾}�6=&��j�3�}�ލ��>���P��/|�>�˟�LMO';�uf����^�,�M��M(,��?	�$	���}89h�H�-IM$0�N���%�o���v�ޅ�O>�ᰋ�}����'}Hvq��1�P�y睋/���Ӿ���hc5^��O#;g�r��]5{J$N+x$�ɡӤLt���k���GM���H��0�j�ql�ƝA���T�̍��9`�Vz�#�7�r��Z���&vΦ���x%N;�R"�POgp�0V�60;��\�b��HgI��!��iu[B�^t�E2zA�R4N�`������x��*�
R�D���g�)'�?yCRwB��=�nմ3�5�����)�mR��+���t9	����ұMxu�)[�hmMnN8M&s�ne�����`ќ8U�J�M�3l��:֑LR�����!�
^PqӚ	�ۑJ�D[)�3X�#���z����y�RvT���� )r]=;�Z���3+cK.�u������5HO�@U��W��}�L��VC��Į]�a���x0�i�M�+u6�3�`�-��+�0����)д���u�u��0��ϓ���&�[dS	��MQ�Z�y(��W�)�%����mq	����y@z��	>t��p��|�7�m'uJ�Lc��[�1��"�M�1k$c5th�O/bv��e�A�5���Ā�*B/��s	E�@vL466�x��A�lnV�[\�C�R�#�T.�f��C��������c�v��r�~�8�.~�嘣Q���3�n�*�*0uh a�Iͳ�Ӱ�k�]E�1<��x��IȬ�3b���Q W��bH���U[��_ģ����t��]�*��G� N}�P�ս���_���~�{:���+��/9�󏾀o��l��t!���<k����}�],a�рƹ�Eǹ��a�3@mm��)�5L�Xz)���������f4�=a�����A���g᪫/��S֡������*>"8sfnA�3٬��^H� A`�z��\S��
Y��O�M��g۩���t����~��-hS��=�S�F�N�f{��j�A�a�ݔ=�N-@e`9�~Ig%+.j�ͳ�,���%�I�+�会-%66�X���|������^������`�)�Q>s6��B�Y�2���_���}��`i�����{u��a*E�y�=��Ycz~��M�n73Xet�lk�IB�!��l��������dK������;M��K{�(\F;�n�N�iۼ0?����֩٠%n^����xz��A��E�ڝ3�q1��t�g�;]N��I�]�N�Z���Yj��}��0ƃ��fA������7GZ�v���J�qb�v���"Si������x���F��y�/l�8�(g��!I�M�BQ8��9��K���#��FN �y��w���B2w>����A�n��cǗ�l��,�mqA�¶E͡��J�1��pǝwK���a+�1p�Qjﾽ��@d��ؓ=3�%7n�o����{�,�i��l�c'g8�b�������l�lNr�Q+��<:���ċ�x��{�0���7��5{����t��N$���d�����V��RA�;��v��D�Az�����#�Y��
O��ـ5�~O��T���ir�Ie&�+ͺE1y��,i�E��L)�77������u�lC��5p��	�j��]خs"�S���ێ3th�M��(�������]{vcq��;�����R����q}�oGf�TD�����D�v�j��þ��Fq�,�������l[�c�l�'�6r��2 ������T	����܆8O[$/Ԉ�N��,c'� >27	Y�5�j٠��+�����1<L�.*۶q+B���^�eh�x�`���d�P�Ƕ8v�>qX��}�|?�<�$��Ѧ,Ja�C�6`�X 9|�8��XE��@�Rg�VY��Dds���	�����F�Ō uv�E�i��c���%�jT/�1e�:_/J_R�'De���[&�-�}_��?�AP�ȶ&�.Mx�����E���d4�_���vj��Cd�4Nt�ۂ�Ř+.q)� �l��b�������}͋�o�[��It@������9ͱͮS�qc'��� �k��h�B6�@��5ȱ� &�U�����d�(�Bp����7�Q*�Q�TL��'5(8�IA�n�-�>�����<{��I(�S�y[�<gB���x��ep~�t.���nx�*��k�������^�V�08R�Q�ss<g�zM��ֲ�6X��������%�U���}G��q�����o�RA���N��Ed�,,�/F*��4��)��� %�C��,��F����.��(���Q�K|��o�6K�z]�\��[�U�hn-��k��w��+.���jz,T��/�
ԡ����f���}�AA2�7�;=k�5�Z}S4���=�5]˧UD�1B���G>�u]�b�."��՟Mk!�ۨ��e��Z�)�`a�e��Vs�A���4셺}�r�х��`k�T�VVVE�9��S�M�y���T�No@��|^]`C[���:t3S�~�8��j��ĝ���@��C� s�d���y>��������K{�*k��fw�y�^_=~󋋘����s�v�PH�4IG��A�>(^���V��_�\ǅ�#�<.ba�*�-�h+x�U�x��VVP�D��Ŋ���m�Bbu�8�]��>s�5��$ �n�`���E`��a��$Lx)�;�z?�|���B��a��ݓ�3~�Dv晭*��ٷy|�j1���/����iH�<of����T!�W���Lij���7��-&�5��}����W6eD���2Σ�m+�NP;�x�1e4X+ҳ~�q�pa8�y(+u�b��9V���:�eٲ���T++k�e�#�"]λ�GH�'�i^y{�g��#�j������:���h\7��?��H����f8���"�2�\ sH�.;9�v�=�$6�=�K.~:N9%�?|���7~�/���;(U-Q���~�����0���S�ig)LO��{�O���$���l�ׅ���8W�s^D��A���T\��\b�KY��x4Z[(0eb1趪���"`t:���_�Y�O���X}��ą�0-�LK��}���#�gџ�K�/kq\<�=d��ܽE�K�V�NǏu�޿�	�����Ϗ*q���ۀ*67Vq��������"��w�B�12@��4Z�R��=
1+1 ���e�w�#����]�qƁ}����~!���uM�&[����S�6�Ųt�z�IFm^U�ؤ���H{-M �hs�-�\=�Pw�e�fl�>��YK1���-Xw~���1�VRg�ߋ���Q��"��Jشr����q��Q�[���޵K6d;wm׮�(|)k�d�ɛI��
5�Q����ff�P���iu1=g��V^��Q����O81�Y$Å�$* ���[�Y ���ܣ'�mԌ�ϲs���5-X8tNv<�0E�qضzE��1ZR��}EP�������`m��~o��{�tL�*<˞�HB#�MM]�v��<@;d�P�'NX$�Pb����d���	S���E���s��`�G�L�i��[Pp�EZ�,��H#��Q*��q�8��=??�ZH{0t����-ŜuO��1`��h|��lI��6�}٭��D�:���g��O���E@�2���s�Z1�K�:7N�I�wu��8e?��6M���K�q뭷�އ�)���g��	_t1�<��7��-��[�RY���ms�kf��P(%F�]��AܟF���l��}�x-�b�>.am�2���"��#.���bձ(�V�P>8�)�Q�:Ͼ�u����ݎg\v�y�ٞ����*������°�nM���{ϲm�MGRE<�(/NKQ����hg�0�?���8x��zyѳ~��Qv�F���\ǽ܃��q=��ϼJ�f#s%��<fv�ڱ ����ЭmnaiyU�e�R�`?a�������a��֏ϠϢ"��i���^o��'����
��w�*�ӡ���uf���`��U�bF��p�Jg�X��qpC��w=����?tt	��5l�-c�����-C^�2I �y��jM�F�et4B��t���W[��v+<u9�t�p�}`�E݋w��v�/>:���-�"�[W�s���������[�!�����̺C�1�����aV���V���Ȇ�S-:�<�;��(n	g���S	=����K��l 	I���U��ۋ�*TN�&kR�<�Y�gx9P���S��iΤ�X$�9.)����lQ��J��C�y�Oao�g͇ݼ����7�mM�ba�t<۵���h�K�\�1�ze\y��ǎ��С9��Y e�f�0SΣ�n	�dS��m��}��������Հ�N�B���»����`���%��|:�x�F3=s�pP;\�ä��F�U�t���أ��O?�z�����[�𶷿_s����x�k��X���@��@�2�V�iJ��3(���	�H��� ��n�����2��`���R�MϸȌWx`S�6�n��H3��b�K2��!qh�f��V��ng�w���?0Y��m��8Im
�{��3��Sjp��j$'"�}����#��C�z���	\ح|���k?>�k���?�5_��Km��~�!�y�ܜ�9�����w�T��ɩ���Q��\q�F��A�i�q�jm+q/�\)�m*�V�ܬm��j�^��/�U��魽�U�L�b�ZC�����
�X��B����<����+��2:Sofjd���P<��Ĵ��zW��T|��sξ�r��C�Li�C'�~�'�T65p�2��N�.�@��\��Z��W[����b�&���@l��^��j��+歝ع��b����Jl�i��uhR�� �ClB��3Ȇ��A�[����ݑ,ӾedA�Z�i�+BP��sW�A! &?V� @�Oh����>�!b��n)�10��@�m�'<����    IDATh�s��BFʅ��<��Z&0Ws�F��&�g�Ye�87g�G*:�l�StC�E�<�0�hg�����^f�tGmD���)3QBd��$�R���c�]���L�`� BL�m��;���K%��1昦C:���(��}�9���p�v��bF��i���	8۬��~�sϱ"�[CƂ6���Џ��1j���v���:f�����ܯ�H8?j�ܿ���
�|��M�}`?���?�;�_��X<�h��"c���A�z�]?qX�?�����q�x���y\��g�s���V���{�(�gU�M��yb�H��M��M�F'Ե��x5���:l�a�	4;��h"ʧ>�IK�vG��=3/ɖKH��N2ƨ�h`c��H?��	|��w�O�vP�^D��W�h�ʠ�.��,�q�}?Foc��<��݇m�;P*M#O�K�f�c(u3��c�V����mfll��	.1ݩ�iː34�la}��[G
�d$�΃.���4!=qb���Q|F̙�U�� �y#:�^�^����SӉl�e2�Uf]��w�
�̨�:J��+��a�X(M�qc}}�Et�`M�AVt6��	���I�-Ϣ�ޭ� H�,����*�^pe��#�K�P��ٿm�j�M��y��phcnp��2�[<@��<l�I�$\��P�b��5鄃�V��JMo���Ĳr��<��W��C=�=�Yh������t�-�[�6	̉׸�\L&6���#�2�;;���*a���+I+�#mv�j��UU�l/zgb����Rat���Gqw`Ywg������N�"vM��7��X�(k,��8o�G\�'c�w�<��Ţ&�����U�L+��Q{΁Q�����8���Gx�ɞ���0� ��4��Z�88�;3�?2��0I��wjD��fK����r��4`vN�!8��S
8z�����_9��ܜ́��ĝ����F�P�0��DI��,���hTEu�
G����<�������?~^x��I\p�:�2>���t���h>e2�����󚔲�Zb�6���4��_X���-�ޟV�&q1J\{��K|_�J0_�!*I��uP�c�����4\Z#�zt��n�.~������3�k�<����4�����ֆIg�9b> v�܋�4���b�m������j��\5�������Qo5P(��Fፉ���ba+l�֖�5�r��	�1�p�v_����oѥf=�]�Lm���e����\N��5�>f,��S��[vsáLQ-�i]3��TA�A�b�l�&A�N��l=�;b�Y�2̥a+	���v<�>�����:��tr���W��,R}�J�&M\��,�4�➕*�
s�'�D�cp	��isցHH�M��"f�`��F�B�����[d��N�������fM^ö9a�/����Y�%Dڱ��'1}+��+���N)d&���V�e�<3¼��߃S�Q�Hb�YM]#1s2�h�e��g&�H�b�e������f,�sیXC�a����˄gd�[���>���DB��n���a|j�]�1��	LB��W����)�uAs�����c;t�箏8s2���
�J�)�SP��Q�|��ȑt?Z���8�(4���H]h�G�c��̲n�����.:�}���
��i�쳟�^�������=x��~ ߽����������)nN�+~�ض�(�;��Dc++*!��Z�ll>��3���-|������&��>\���X:z��v4�5l۶���u�{n��G�?߸��O���-L�8i�K��5nIY{D�F�ǰ��P��[?���(SHw��%#���Z��`��M�[�3�CVٹ����$5_;ȣ��z�C����s��Χ��\��v>�A���|��V}E�TO�k���7�gfj=��:�Ә���"�v3��,���	��n,'{!������5y�1{`&�`IN2'�� �8���U����-��l�H�p'H��j5Ӱ3Rٿ ��#/;3,���ahK�34!� ��4�;Ҿe�'W��V@eЉ�H���P]��aoJ]��L�A'5�����n�f����NF�*Δ��PH��k`����$�O���]�d�8�@Mtf�!Kf@��w�q�u�Ns� �g��������>�U�UA�l����d։
�	k�A��q�.�J��ꜲH��`��\t.܊�r�߷���=,�}&0\L�94�p�̊+�p��l���8�-w^2�eםC��x�-:������pȘ�|a���E@�����8�d�M�0q6wPt��2�g���Ți4�ZX���P�Mb�P���o��G���~lJ�v��j�fv��ͬ�=�TB�\Z�v�{Q+i�Dt�Ja�Z�m��}T7�����A�}����\{�ɲ~�/���^����x���?�}�x��'�}�^��W��k}����Q�g�q�#��YB�`��}������%.<���ȧ7�B��C�;~����V&{�(����|�>��oV�D�4"���$���h�s��s.<��G����Û��t��Q�ѡ����V� DF�)&\PC݂^��3L�����e���;�>�O~�0��9��-��ӈ���F�UO��L���~��a��W�΢4ţ���e�Z[X���z�����P���uA�(t8nm�U���M���7��8�	&-ᨼ��������!�|�]��7w��v8�h�`w�-�Z�(SX����#��F"˼Y<�µ�?@���DQ��N?5[3��<��<�y�2l7�����.�E�.5i�A�ޱ�=S.]*�1�!���#*,R����E]�BV�3q��,���0e:��Z#�SA�$ ��HYӂ�6a����"d��R��c��1i�0q(�A;llF4�̓��aMf��� ��=���;��\�1K8�m���v��(,��v5�0@sE�e2^PBv΅7p�9�J劂!�v`y�5�>NJe�Mhd(���i�3���!z�)g�g�e�������GJBe�sK.tB��&K�s�y��j���L�����<�$1Q�m�&�1�a_�ۛ���������5�R��!�Q��*��UW��������������<����J�sN��|��6�_~�K��������=���He��+}�|�m�\Ȩ80��������I�NK�QJ�m�(��-����m�x���;۷�j���|���Ͽ��h�(F��!�~�fք1ҨՎbf�4tH4�^t6���K�od]O,���dp�fXKx�v��HTe�MYx:��-�v;�oG7�h�-q��ъ�]��h�����%��n*#���Oӊ+�n���1l�(�3Q���6LY�����<U�G6J|U���(i��%b;t����*���iVWsl�g�l�l2G�A�.�j�ɤШ� U�&��N�ݘ8�=��D��[ē�A̓�Y���H+#~NL.��B<X��:�>���5A.�1��$X�����.��`��Wـ!5���۲�#(.��ɥ�:��W�j�g�t�[B��%:�ټΣE}�`]�AY�l�Q7�6�Cl_�NJu����@�(���	���Ý�v`ԓI����L�]�nS{�n1BQ�M+��ǿ��1��Y̤^���#4�`n����=4���`�/wl��z��q���ِ��b��$"�M(L�IR�k�uQM�V:ݑ�bJ8��%$_��Oڿ��<�CA[(	7˒�D.��vsI������ �pȭ��A��y'=$�����9<R+6O`��m�9`#ì�|��ES;+6��/�5*�ddx���s���]��^�?9_������?�����o��mz�t�c���
��A�-����>֖�{��\rqٴ=z@T_բ����E�CrT(f�ͧ%�u�i#�-'�u�|ԗɦ*�XC���aCN�>�4�ƴ�jؽ;�[��"�{޸c�&
�UǬ�G��fhC�D�c�#��c�ufI�ԃn��"��:�0�Π^�����@t��n�5����}���\���`�V��;뒏,.�N�v��A��Q�;������� cⱶB0�h�j�n��<85�yj�����^���-Ӡ�>/�<�.��N��8.X��[��5�6�4�c����P��*��3f��X��u������':���	��e�.$3W�H|���J#��:[��#��Lj���l�@��z��R1�%�!f�%����8;�dY))2��UÀ�n/����Aō4-��w�\p�R�B����!_#�ѱT�O"���b,!
�mL��
�Ҩ0���@Ѹ�d���l���;�ߧE�N�p��	���7�������]U!�!��"�b�kܳ�ѓ���-�=�Qa��5���3�@�$���X}&���">��{�SI ��H���5��a�*������zj�%����kR{�b9�bl���?���D�j�1LĤ��{��(����m��+����
��Dڄ�;Y��MF
�Oޅ���W�/گ��vw�|�	�P&��pc�m��k��i4�=�����Ӯ�g;h7ְ��^�������-����66ĲY]^��-g���!���D�@�@�`	�w�}w.����1=t�n؇^!�Nj ���;�B>ΡѲ�fu^��_z�s�O(���e�
dv�<�M��Z��<j�>
�[|�o���&T����geg1�ͣ�ɠ�n"�����t�zQO�M�!�X�>{��=�x�$R;����T̲F���j�aA��]�+&�C�9��}�&����2u)����T�LvP�f�T��?Fr)g�#ޥ��[��=��X.9��W�����%'��I��9��>, p�pr0�\����:6�� ,�"�$Nh��N� �r�ﬔKʰuĶ������1�
��~����z���?��-�b�x��)Ժ���q1�Ow�ٻ�/L �d�T֥��p-+
�vR��2 9�B�aV�⠧�0E���r�k�Al>��G����M��	IA�U���'R���.u���L{�YF-�~l�b��gQ��njhq0�W:0�:��0'vg��)Z�NS�wҡ����;r����:�ӄ�R��ZcИ��$�\��O�K2Lʰ�І(����SĕV��X7��?���4�m1OX��#� mΈ��u�u�������i�d	Z����a�����&>���I,��.�o����o���6�t)G� >��o����z��rq�`ZQgi,���1앰�!��ލ��C���m&�T]�[��%b�(h�=����X��#�y<��U9E;��e+I`�N�3�G�������w�E��U/�7�t'����4���X3=eu���"kUҢ-h����/ݮ]\�m:��C�ؘ��Q�Ċ�ϼ�GC���&E��aRŹy�d"�i��H��E�������ٵ����gv�1؃A���Y�t�l��m0��{I�r�1Cr^+��R�k6emd�=�]fQ����p��`�n�3k�1��5Tʭxf�݇d�~�m�QJf�f^J��#��ˊK��<goرm=���g�j�?�z@�4O}��,25�N����EJٺ�i�c&���%���2��`�Y����L�����"	��g>�g@�� "�ʔ�4�ʨ	��GY>;T��(G��22��,�#Ưݖ++�]��ЙFl϶x����!�%n@n�5$�}^���-X\��@>?�3/�>oG*�]�j��c�k�%4�u%:��&k<2�]�Y�)��Q*��]�.��Q& a&T�:(^O��"A�b�n/VCa �uX'�Λ��jw���_�
�
�I���12 �;q�i>R��;��N�b�:��W$�N�'���:��!(� �
0�ks�ʛ6����eQ̦�rdU?j5��Ͻ�fw�/_�]��՛��O��M���/��q_���h5���nΰ�];L�n�9���cs1��ތŅ8���XY=���ka��v�.#��	I�J�a�c���1n�����7��#��hD���2�9%�`$��f�No8`gf��$߾�w��Uػ����x��G1���<�ع=���6wn��� _�Ɲ�>��k�)��C&SA�oJ���t�)������-��~+�:Z�&�b�r;�l0(��N�"4T)}�X
.nN�����G#�F���@��.l�#4Gt����,�2x(2{rL�7��i�wzu��A��b٢.��=���vO�A:e�°�"bEL����D57�|�ƪV�a�,���:?SLoI��I�].�r1��	q��lD���2� �d���¬�Dg�z#n��Ӽw*��V[�����bxX�G���6����k3�-��k��00$e���0F��Z2��L�C3]�U ��&Nb�-���n�x�D��VB#衣��� 
Z�vs=]C�g��s�v��!�E��-�޵ӄ5������Ylp?����Ԃ[��(;���n�T�%��D؁F�z3m�y>�o&��Z(���A�T,����!�[�`�����nm�,_�-.��n��Mdۡ�G��%Lf�����B�	��@�7b��� %Z�(�	�0�kҰ�Ŀ�r��
�I ��XV4,���a�ӭ�2N߷�>���}2��Z��o�+�2/�_������8��w��~�Cx�_��|�di� �����Aw��1Legp������ǥ��v�L�i�07+��u��R��Xu�<_�m���6�ggp˷�C����r�9�6N�ջ��L��0���$����2��^��q��2�%�5?r�*ǫh�ų�y6n��O�Ա:����y`�QA������z=}s��Dvj��O�<{�#��7��Mʍ6ju,?���.��"}@1afʂ.WӍ5b`d6��^J�v��m���	�fq~^�?u�䋱g��'+����I133G�s��,��`~z333��`Ѯ�"M�)�HX�0���5��8��&�,Y�@O	35`�� ��-B7l�I��q����ٌmb�&��lgٮ����Q�� �<i���Q*�`�b�N�ȼ����j�k�!<,�tk2nIU��'k�u4�$L3ƫi#�K��Y����L���Q'�����fj�O����6�����{��͒�Ґ�M�LXm�;'.Z
8�(uP#�)E�(F&�9uݴCF�Ie��n��������(vp���h,/k'NSL2G�[hQcF��[��B�s�qGq'���U��Ʈ����x���^�܌�G�8;wcg}��v�EZ%z�u��9�9'���ƭ��7��a�+��w�*���'��Bা	+i�H�!P=����BF�m�.&;�f�\^::T�z[
�o���⳷)`k�o,�5?��R���tpli{NٍO|���=.�t�w�m�:�31��[Z(��_|.�z����m�,/��5&��ܴ	ҩ�[�i#N������ ��(�ը��_��f���c%��o��uh��r�rw�e#"=g��~߶u���`Ϟ�Xjcϡ8�V�vmK�8��3��t�t�l�^��<����O{�8���<�+�%�1L;��ۡ�R<��>��]�p��X�����1�I�'6�b�*�vyyeݷ\V؋V����) �'��w:֘���@�m��m��]�*@�ܱ��}���l�s���F��]�#ڍqG���E�_�I��f�e����$x)JF3��T��	�b���%�)M눓���k�	�D�9t��:�>�[������>gh�qB��I���>*/�u�e��0�͓h�ڨ����(抨��*�p;��l�r3�K�\z��]��s1*-$�|�@΅����K�ςqƠ3.d������5F�����4��"�ʫG@���%p���	Pۣ=����/�RO@�U+��
jʓN��mA��K��mu�1M5tB�p�Lt>7�X��}����M�g5�5A+%�����*��C�W��Z�Z�~u�����"�≻�㒍Z��A`C��!Z�CS�t߱X6�s�$��?ؒ�n{ǣ=�`�fi~�T��<�E��5!�:���J��Y�oV%Ey�    IDATA������4�Rb��s�=��)��uR�px<�x��n��{�wnt��d�S*L�X^z���[���E+�Uז�t�!O��g�+RbGH��g]�X'#��D�[»�kj��"MS��Lυ����t0��o ϿRk`�{&WF/UCvM��h���R�H�����0=�UG��e�m/j�#�&]��Giv�g�o��f��G~��a��E�~ک�����������6%�C�9��ǆ�z�%��V�h1�۶ϩe���V�&�A�MjۗkR�sW����'�����<�}X����Z����d���٘��3��Jo[�NAs�a��c�C���'c3Q	�xf�,��<!go�
�}h���n��%6H*}*=���Ѹ2�\�Tv�V����Yfo����l⫑N.&��&�{��kdTkt�:��x��Ezh��=�ﱈ�@~�$i��,��R��[~g�0���<�kL�������b�\�����9�.�h*0�e����{7�U�?�]|l���ÄPd�]BW�3O�\9�Db[|�%�Y�H�h��L��A=���V� �%���Pv�1bs�#2q\�`��n�!-�N�L�MoI-���!�yOUL#Dŝ�u5�@Dc`��XoA(>��{X�6���H�m��t��yF6N���Xw��8��~o��"����j�8^��p���b���D���οt��DFX^���&۽g��8SD&;Bw��l��+^u*^��gY�>?D���N�����7IS��<YA9t�bC�������KH��g+�Ȱ�\�%�`�.�9��C�,Nj!t��\w�t���l	�a
�^�aQvy��ǕEIhs��\ ��$m6�QVc?=P�+��׳AS�方=�s���-�Q,b�g`��ff�%������Gʒن]@�j^U�`�\o4A'����̓�,0��e�	+�ub�<y�I�X�Ƕ�yĹb2���S��6aT�� ��$�)G�qƠ��LG�1=˘U���X�<,ñ"�Y�r���a�x��F��&kҨ@Ɖ���P��2Y�9a{a*�l�L�gV���A2yy��wP�ܞ���<e��s�"�'�������.H�l�=��g�*�j{�!�h3�&��\if�:P��+�xn�-1s�h�%��y�F���D���׹֝v*eh���닐	�'t6q���6��w;�Px;Su#z,}kQ���="�b�X�v2hZ`G���V��g���e�aQCAE[�|����!�7K�d�A���l�$�D&�׃�L�0�r!��;}2{W׮$�� �3�yhl{>V����5ct�i$���Xszc�Z=��a�N2W!+��OB���t:�_������C�
�q����]����[��!~������C�"��ۯ��~�8���x����r�j��ȧ��3U�#�h�ع�v��.#�&h���&�jӊ�����MWe�x?n��ݨ#�/!�/ Om=�����܃�.�k�7a�c�6�^�����vj���Y�4Jӈ502p�YfH�Wp�"�II�!&���q��肗^?*��u�8x���ol`nv�^�t������t�`f]�����i���z���,���2U�]p��a�WM\�ۗpHtJ<锤HI=:��Sڎw�]��L#� ��#�b:X�U�&v&�Cb�x&cM&l��p̾|���dEް��<c\i���I:\����`�w9Q�C���Z��Q��L�0q��VZ{.q�Pr�H'F��4z�ru�LT����X;���ɑe��a�e�kR��Y��)=�&�
�������U�dfo�a�4h�˓F�V�L�¤s�>ʲUTQ��U�P�$W��=_[x��e��LG1/�avͪi�q�
�I˔V��&T�����6���ү��ƮÁi5���Z�v��Z�M����t�)~Xq�;Js�7&]�5�:㤈��u�-f�͆qlu�|l>M�m�ڽN��oHl7a�x.�<���������ҫ��k�>7�g>�n2F1U^����moye�@��G㻷܅��&^|�K��{�>�Tj�31��i)}�n��F�a\~�~��;��m��-D��`��Ĳl��y?�>55������w��k�Wff����c�N���:� ��7}#�y����d>��Vi�}�ۂ�3�<J���C��jgd�M��u���*�?=t���/�q���n'�Gu}�aǎ���]����?���U��i�:�Y�G"���yĕ��9��3�(�Ʌ1�BÜ���j���� �">�Q'�WQ�C���4f����y~�X�gi6�'�O�I�FJ�g�3��� Ek���vi׉A�V'��d�̏p�&{��|9�BFm�,|� '���P�̈́d�E�߉b�[e��u^�w5�A�c�d�$����(�R����i[=���;��>+"���V@�|�[v*(�uv	�z�Zcƫ���I�e�a��`���-��q�DAQ��xAT+8�٪]�X�Y�Do-�ő-P	<�E��!�+ zC�=�z"!�mυu܁^'E91AX\�"Cg�����c�;���`�f�':瞬�zI�DCj~H(.�^���A��zK�A�`DF"�w������B�
��x���a�V#G�S±�{��K/���i��ê?��ϡC}�t��˿����?���� ~��᪟�J�9|�8Rqq�ھ}U�F$5D����W`���%0A,�0�5���s�.��m��5�ry�eť��A���?�(���lq��4�M{m!MR�XH&�~������7��19�>		1�m#���9�	q1�wjws}��
H�ڠ�t=9r�(�u����D2f�L	�yacuEM5T�*A�1�m�n[��2�<�-o�1�>�
&�Ww���0�4
L�lUB�*�9q_PCPܳ�M<��� �B�=D�;����is�r m�ՙ
7��e���v�\��R�R��͵g���x�)�Op�08U�$Gֽ��V�6<a`[@1��D����L2y�< 2h���A�A����	�u��e�!K�N)-���t�h�x�iDa҆���!�
��J���s���,	U{���:���W��]�8p'P~��q�]�I�=A?�����F���r�3
ٵa�b��0YT%?y^�IgK�-���Y�0�/l�s�̯��։)D2|i�R�i���c������-�¢�Q�E_�=�lmr���acsC�I.c�Dc�0`n�:M�1���E[���,D��n�ȌE��50���Cҹ$�!~/�n�ﲷsg6�m1��y/:�z�5�(Qr������������^��׾�����}���H�8x�At�M�N��h���e�@�QM���۲�F��چ��=���|շ6P�̢�>����س?�T�����U?��a]]E&_T����*�Hr���]s�c����V��	!��G�]���4�,�q�
�V���D=��8��⵩Q3�]���C���-�>к-BN}E(O��5����v�X��@̊+�+��{�D��wh�x� g�{>P�Ѡ �Й"�KM̩
�I��iaH�X����%�mE��&d0)~��1'����c[���cg��=�*�ξp�=���a�	;w8n�زn����a8�5����-���:[�y��tHqJe�cH��1G�0����I�I6�0[�������[�
ߩ��#��#�gl!���5Ix±~}��R����Ȃf��?9�<X��2�ۭ	���>OX<tS|Ga��wN�W#ǚd\=�m��d��ЌYi���r,��g���Y�4Y�9�E�M��0����(~�=Q�ċ�2��@����%�>&:l �n[�L�@��c���1�ܸ�4ʥ
�z�t4d-M���EC$1��物*&��:��V�6u���A�\{[|�1FC즏E���҇�?����m�;H���SX[9�7��gp�˟���s�Ԩ�k��l!����3� �ccs毽��'�i��A�vbx~�{�~	�L�w�3��/z������\av6R�����ЃObn���e��}�����l%�`��|����y�{%=#6��]�J
&�Z�X��o	1.�[��3����x����3�J��2H�c�b2�r#��=i��
Ȣ���W�8�2��Z��4�c���Jp[6R��M,(�7���\��]dL��ޢ�&3l�*ඓ����Y����T�b�m��efV�A����g��l	2[i��C_��%7��eƊ�@4�U8�L��3HQ�����6u�Ԅ:`2�m����j29���E��D�7�Ȭ'1�kÌQ�k{��p��s��:�0Ȥ�h�P�7�����"d�f���}RT3���k 	���Cf�ζ�����8�ψ+�t]T�2�7+jY�F��8�ylH���a<m�+��Ķ�!�N��d����]��pj�֏��
�l��.걂$�����T�o3�#|��c^��mo n���*���
��� ��uolnbaβG3i��fo%�>S��'Vg�y����R�����vj�!�]����[U9��yLMQRߞ;��}H�d5@�쟺�?�L��Ti�k�i�ư�X��#����j<���Q��c炅�Y�!��U���߄z�(��0�1o�,��؟��U;��.�z�l�]��j�_~.V�7p����G���3���hh�w��B2�Z͆���<�sshw�¾�y�<�
�¡�
�%�k�x���x|'�v؅��)،R�`��>�0Nz���o����V]�
)r�����~�+4ul��2�TS��)"}��/�t����"m)���*mD�5� �s�X��m�u1z�$yH���>�b[�_�n�}����!�؂��´��P�mf���r�1-zd�M��[2�<k��pɃ�
3V�y�LCo�؂�m��(��B��|X�
�_��V�m�,�h����&���^�=��	1s5`Xᐷ_{\B)�
e!��EHV2�AQ��E1m�qX���4T@s�a�5Z������:�a�k<0����jc�������ߎ��t�}����-�����P\�m�LѲ�������Hmv/��	1)��𦕰Bp�	��x�٪ډˬ
GP������;��UVx�owة�q�p�g�$s�`̃��e��]�X^��w�\����F���y
�L�U�x�>��ٙ	~$���tE�/��ڒ�p'!x|
a*�g�T1sG��ۊ�>+s�5n�n!�//=����q�����M�G�����O4�{`�y� <�D�����?�R����8��A.]P�ܲZ��E��G��E��W��
|�K�a��m���9�رø�:��Ycg�ڎ��<Fy�m��9�w<��[-)Ɏ'n3pso�cF�eӛf����&�#�g��SC:�S������6�H���0䂟����F �d�z�_uT9%����Q�����Zy�j`?���0{	|�i��1ư3\c�KN���A?��oL�A�*��D���
<�E@r`h���l҄�Ǉ�"���S��ώ�͛,>*x;jb-�&줬]���.%�`sO�r`�5�p�{�2� ���
z��9U�$�âX�t�Ř����G��A@�:�|M�4l���H�6d��'�n�p���tc��(�U�p❺�r=�F&\�qs �;�	a9��u�)%AOY5?˸�Z|\�[BaW��?Y�[X��l̀B�A�f��lAR f�y"tm�O�IK��,kB4�N����ŀ�J�|�!�Q��x5Ϣ;0
,��?�:�-,�څs���|ϸ��D-�\�k��~��?@����Z�|�y8k���F��_����U5�#G�+��i�d|M�NaqnVA[F$��N��r�AQ����@�1X8�U����X�f��Z�,6���h����fL�����)|�[������e?{����=����o��Ͽڸ�3�����8|��|�����R)3/lX��A��t[Ut�����֫�[G6�F6SD��A����_}����0����J��2ԭ-��~���#�.��M�Y�rm��Hsc�̦�S�3��t!5�:|y0ـcG��Q~i��i8�ȑ����j6�J�}1�W����p�d�*kـ�����\�\���":ТuSl�݄&�2���2MQ����E��At���3(;{�6gڠn���>J�:���U���pMca�^|�d*�1�J���m�l��Nv$<��A��&P%�n�%.��fl߾���d��A��c�6�V���Avb}�L��<��bƏ�dM��m*�Q��&�]{$=!�2�Qd�^h�+QLC�&�1l��t1rk��Q%���(�I���R�G�F1
�VA���u��N�o�6��`�9��i�gyXj0z����L��~i�X<�$Ayoh�l!$�˰|e���/�:<��kQlA*������ ����ĳ�O�K�j!v��Eek�&��;�������,S��5ȯ��j9�H�$����L��s�=j�llbv��r���.�H?S"4�"V�=�F��GO>�����g�J	�33�f�.��pK���?j��k��	�GJ��94#�@�#�( �� 8���G���^��g_q.���2�?}
'�7��|���r�t�C(w .Mam�Q�{�;��hAϽ�.�1l��n#�b<��(�ڨF�{+�4�.΅��\B�������d�G��>u*��~�L^���3E*cC͠���	X��NX��Ca]�! ��T�����(�f��A\�R�y>~�V	۶ȍ�T!�yr'�F��SOIѹ/��H�״��p�A�j�Za�Y������슟ˮ�d��\3#'��n,*V�u<G^��b!&�x���������'�6�H��@=U��A�q�P5��;���7	�=��Y�D���F�������Ir!c��G�=�		��&,���4JD�.�L�4^�}�MX��}f�NUS����
P�u.c^�~.����pa��GM�B�J(�ɒ�~N����{I/sް�8�l�Ť#������|S��=P���z�y�$�d�A'�"ӊu��,8�$r�OdS�Ԫ��W��P	O�z$܉P�O�F�S�����D��,�"Pnѥ]�O8e���L����6g����hp� }b��IQ�
����*��1�'�A+�e���*p��8/~��nu�`�qS�����#ld�EnmsS�Q<�q�y(����J͏J���s��1�/|���q��]8����w.6�:���8�&�������w����e��jU�|���E�k54j�b��]�_����oz�{�t|���^LM�4A6�Ǳ�ǐs��Te�4�9gzцޗ�I�Kc�&/:B��8d�Г�τ�N2-z���k;={l:�He�{��Tʀ�E�.Q�5�IK}ߕ!9�hF�1ض�9�㑳ۂ2�Gw%�̕�f�� �i��?�P2pF]�2t�C�� �G9I�`!�U7J����c�hq��$Y��"�6Wa�80����Jڶ�zR��&��%}�}���!��	Vm�߁�z�X$
N�
b�}ϺX%wQ��%ʀ�ه��)���j�qf����Q��~�s7� �Ia�K�A)����9Y[��*̘��&�M
�l/W��5�p���4��l�U�Dɲ�����4
i36�u����R�i^*a�54{�q���.J�e��2�� �aB`Z@��K�P��U�oƝ�FD7<Xa�N9k�]���[qT>����#ӲEU�4#������k�2A �>7t�2hSwD�T�ef# +�y�|L�4+,_5YsZ����3�:�5g� ��;H�{�}���4mr��(cbE�s�[l�'���C�<��O�+}������"ʹ�QE�[�G1�_V�sec{v�Htꙑs2!	R�ܡ��ɧa��yeٛ[(W�|�A���&-ӂ�ɐH2x|M�τH�)��F�;m !@޿�(뛧3���baa�k���i�,    IDATN1J���݂Rы���r�7���UŶm�T��.�;�>��Gl��Q��JYbj��dS�EhHYV�h��x��}�reH��n�ƠHlEs(�D'��Ս�'�/���Ȃ!-�;	p��]��v�:�}/��x��2o�&s�"��fX$�e]$�D]s��#<�{�Ĝej��VxR�&U�"8��j����$�m�qq۪�����OMA��"��^X�*Mۺ�A��f��p�Y�����-��I��F{OȰ9��&����n�hhN����U��t��癑������s%�fuƹ�!'���U�e�v�1S�[�Y\d�X�v��%#n�I�O���%�����+�$���;N�݌�O�S�
�b� �~6��_��l׳�^�<㙧�'9!�����B@D���������T{��j{Y�V;�D�NT-*Eq D�$$���'g>�����w����<�^���u�|�;<�}�{�k��V�c�M�V�d8�H�*$[�iA$�6����[�8�Nʰm�"Ӧ�BѺ 	q��2�J��ƅV d�嵊��N(n�Fc�m����zw�Ij"☻w�w\�.��S��l�>�K�v4r�d�&�]�yC�vޟ����kk
����z��nE�s1��T��6K5Nn��((8=���j*.O0�cgw�rQ]�ܭ���|-w�1g����)&X�=�L����c��x���\�u+�쮣Tn
��d����M"�����au����v��t��\y��Q���%w�����)y�4/�=XC9WCK���3B��R*Ug���Wj�".չ@��QD�V�t�dF�P�Y�P���Ϣ�
�ク����X2(��u4�Y&y,��|nƺ=	�ʸ%o0���#���@�U�I�^���0�TjPj5LC��&:�,py�NAN����P4�;����)S
9
̌T�0w��m�`NZ�v�rz3��VG*8�Cܜ]U��V0r�T11hf���-؛�E��0���:�8��T�(����:�P|��m�E��s[k&e]i�F�s$�/r��@��Z^
�p�|�a�!>d�=N3���M<�����H5^?3�)��</b�#k�vx �;Ӆ-]����q�8d6Zv�5$k�VP&�|��S����ٳ��b�On�4�l�Ǹb[)ۂ�3B0�Lvn�h!��X�m�d5�	��� "�C=9�52x��huC�����>�����9]4��BS��LD{�ě9FX�Q�ww�`�n�#I�Jն�M)�N6�8��o�T
-�;c����Sf��`���5�1k���yFH���G��صZ��A}�� �%���m���C�]�J=�ȳWߗ�2�ª[�X@n;��E����lĢ�3_��m�F�֊s�"�C���"Ř��`�`�l�
�A��Av=��Fb��8Q��sv^�z����X�N;(�br��6W6�=�2����p�\lL~bl��Sc>���	f�l�\ɺ�y��t��b�{�l�bBP�`6�!�ҷ��e��*��di�&@��htL�,�m<�k���zG^�6���R�N�K�XI
1��Rǻ�b�td(x#��P�6�5CxaR�-�a��m����:WV��j{�:��>�z؀��b��{MϚ��[���+�O5O��lb�=�k�͗a�x�51�D�ϱQb���P���0kB��&����H�jC�7�+�V����O�������0�k�H��*�2"��@�<��'�U��"t�Ń�3�.r�`,��Y�9J�E.����l�N�z��6YJr�>_�H���/ ��F�2�h��-�4��'�ⷘ���ߟը��I�0U�l�A[�z.'��-��Wg��!�����>��D��l�f�$Ӑ�6���b�y��Y�:g+��KDhB!�"����I��O����`�v��߶��<��"�.Ⱦ}�Z�]�"v���Z1W�K�(�������/!7��Q�Z�f}��-) 2�s�ݤ�k�� [e�2����)�)`2�ۢ��n�2Z�F�:&][��<��w����2��`���2���S'�5T��T���T�Z0ܹ�F�"%��k���$f0g�X����%p�J
@8a�[����}����@�mg��y���#P��PD�;B������zX�eh�"b�l��#i]u���D�Uq�·Hw�Dt'���o�Օ#�^�[�г[�kl�>�]�f��Ci�Z�MPE�:�!Zn�-�c��yα�˵./�8b�&�P:"�"_`��R�b(</j�����
��V�+N����j²����l�p������b�XҸ�G82:X��u%�Gi�Q����W��&��jMZ�h��3<�<8��#L�L�[X[���Ɨ4��@�H������^D�NaR�e���a"��LFE0��	��L7����yj]p��{C�����އħ�����.�8#m��xS���23Q[����,uW�ܩ)�}	� ��N�z�
��s��
dj��w���ӌ�v;\�h,�C=r&��uDv�F6�Z;g���Ιu��ղע���c���)�����k
�Ŵ��'���B=�<G�r6���Р7F�A�	.�f��k��JV�����Y�2�u�4�A}:1��֭W�������f}}9����v����;𪯱"�g?����8~�6���s7����s���={�;�:�U�?��T������7��$^R{��GG��4c�%:�j��kkF�E��F(�!��#̼#=_m��b�������aR��6W����<6$bS/
M�>��3��u�qe7�3<nU��N/m�f\Qݹfd+�!!b�� ���e6�B�[xJ��V>�B��`����E2X�&~hd���9�KIBB<�l!w�L�,O�G{%3��6M���~��:}����&�g���P�
���b�1�N���5%2rL?f�������K�6'�@y�	����ܜy���u���9�Z��Ƌ��L�ڻS,>�3�+![��DJ�s���(���Ke`�����B�47�똣��MXvQ[4f��4��	�
�p!2�ˡ��zf��\l-H��H�WI}P�LF1T�ޏ��+�f3r��a(O(#R\�bo�6�_����^��.�p��q4�`(F�a��RU���Ք�� h�S���Ň����F^�����Ќa�);ۤH+z��b�[F�*���Pad<5���d�nӣ�CQ���C��Hs�j[�.H�m˔6�����;�"={�\��Hӏ��;�������b���X,L�X*��#Q�>�x���^`������7���"J����R+a����DL�|����l����w�a`��#̉�'���<�q��l���e�%̦\��:/�s�_&�����ߙ�m�
e�<d6�L�[Ju"�`����x���edxX���X(7�V(A��fFY�S����՞��(����j��vgЋ�{l
`�N� ��ZM>T;s�Ws���
����.�)��<j9����f��Q���q"�$ZC/I2
8�#d�q�樜@	��:��1�^4�H_�X����c�D*)�6%j$�ǛS��%U�jļh�F������2��~RD2�E/2�|����]<@{��VY�7�xO��u����8
@,"#L<�|�7w1	��8e�x�ɯ:�հ<�4�)�b�b��o8�ʵ��7�ia���.lU���1%�k��졮Q�D����l�k�.\p/�m�)<�1 q�̠�%.63yӡ0�/?/�B�Ϥ4��MB��E=�}��8{��q/u��D�9aK\��q�.��ں�E��~_ىj��Z��A�*���h�Sv�_��ŵu�ņ	����yoi b?1��܌^�%t�=�H��q��~z����W�ě���F�+����[Ke<w��`�c�Mn��'~>lI���!��ϗUw�!c��$�y]���+�M��z8�����MP�7���f��U?ΐ'=�M��'����e��=j���c�;���2c���k�43��M�@>�é���!�Zt9��"Ɔ�pfy�1]k�d5U!.>ŀ�j��A��CTD�l��2�ڹRE�n����d�T�u	%�0m�,MNNj�N��8�����& ����e�&�d"��N�T+ҟ��h6��Ƚ&��g�3�'���~<�(��0N�|(Y$ӽ�^@��B�L�gI3�}�PB��%����D�����O���M֮Iz#�$Y�*
d����}�Xi�Z�]�o�\{�kpU`=І�2�L�Le�6���%���b�X|"�G��J��qXK`S�0��{79�(�<hN�����҉��?��<���-�M��)�d�ZP�R+�ȺL��-�.��A��$�H�]�S.
$�|&�:
\R�� >���F�ˣ���gxб�����:��Y�:�q�Q�J�V���T�qH����/v�,����ư�RrN��t�2�<� �h��#*��,��{}�Y�]���n��(^���XZ.`c����$V�g�2���c��#	7z4Rz_|�,~�}�]��3�t�XX�#�L[�`������̒ٗ�)kkQ��n���	���F�Bу���l>�7�s_�΢z1��<Wq�7�ڼ� ��IBWM!X�{f�$;Y:���3Ȑure�Y�;'SA���x�-L�}L�0�*2�7�EWj6*FAt��Z#�)Z&���k��u�]��#ov��2�kz��mغ�lrv�ZL�P�����R_��~\�����k�V1}o����Ҵo�Ҵӿg�.8+�[�Af�����:�D8�вR��R�#1�;��6Z"�l٤3��8bR^QX��6 =g��J���uΨȒK8�J��Nv$��X$R����`�%:uO�Z��)f�B[�*���>������!�݋�=�f+;�ԥ��hc��D&l
2	T`P!���0X�f���'����,1x��60S`Bv�l���t�
+֙t��ٓ���U��)2prя�P��{�����[]��{��g��x��<�t�L�>1�Ț���Z����R�٨/�ਕ+R��\��l�RSr�x��]��h���LRv�'C�>��Ǎ��ś�y%N�\;�5?�S��һ�.a}g�֊��ZZ�h�Sl(�,����O�¥M���q����6Po�Lm�!#m����c�p���>�H��\�&���;	��x�lY��@�����=��8�̤���o|�<���1�[����s�RG@(�dBMn����P�Vj��&��`��.�ص��K77���6��K��F�h��?�������K�b��|؆۬Z�W�U�H�z����%�C�x��A6�čc��U�X�(v�MX���Yn����l��渂Ml�#4jUu�6�j�5j�R���.\��.�X^}�a0x31�+5�����j�)h����Q�J���t޵��N�\Z�OHs�q>��CŽ���4�+�0��f��f��[vP*�ъ�1��h&ӎB��A��>�,q�=��o/��Ƅ���(�jr#_��_�0��s�����)����5Y���y(5y�fEW5Ll��;J�è3��6�4�I�G��C�[����o���լ1�Bi,-B��G��_07v�A��Q�W���kv�5�{���SqLo��-}1��A)��׏$Ɋ�љ���ޗͮl�	��?%a�ص��Ŧ��x�Ţkn���v��Ϟ�dn"g��j���Qޏ|�E�*�	�)����}%{��9-��~\<�Tbv��r�Q�/�F���ރ���9ʯ�Rȣ�~�?������r%kw/W�}�QeX�
��q�*���
�t�X�����/(�L��r�c:'�Z�h�F����`H�Kc���o�{]t"B���Q�vгF����6�+M�f1�N�J��@F�$;�QT2O: �t鲌�/�����k����}��ޠ�U��4�;�β�0'YVT;�s�1s���$0�Y�S1��f���G���)�Z�l���0(��VَW���V %6 l�m�֬biߢ��Z�-5����k�����\��1Ԯ{��%��[$�Uuuv2m�C5�.�Fs%�b��� �8���J���'a�$�;�F�V��n�\x�զ��>��8F|�e]�d�k��+��β�W�č9����=b���* {L������Z�sX�e�	X�\l�\ˀļԙou���i�-��[YcFX �L2��)f��b2CSD�ee�/{�=2���sP���g��b���E�f?�
y�BR�~ f�`�=c:7q��JQ]}Z(��#���?n�a0�������#��˧0蓱���,|�]8a��ٜqݪ��3<Zc�0Ǽ�f��n����s�}"Å�J�ψ;���o�s��c�4A��o��W�}���eX����a{S�/_|�i�rS�]�X$�o� �ƾ��b��v��FК�����������X�f�ȩ�ֱ��നB+2N
y�Y�a$.�W�jCt�T�[@/W���ݲBs��#�A�19Ek���{�~k>�x�e�E���#�.�r���p�hU6������6M��ɧ��{ٍT�U�v��D�y�ۗ���EI�N�^����e��n��҂��N�N��t��D�l [� �'A��{Ԝw��٧ڴ����Lm�6���q޴!z�+u��[���͆v[;�@�Qf"���;8� O�8�C`64~'U��pG�D�e��\[��UD�����^��s�U���v�N���T�F� m�D-��WCɥ%��ֲs�-8�����5%�5Wc�|��3�*��U�~=8_�Q�g�M��D���������� C>�*�����
�^�T��`w����e�v��D{$�����2I�+��L��em�ji�	�zm��(�t���3hy#u71B�I�_�N���)��蚣B�w�r�Kw�vE�1�Pc1�O��g�Ƙ�ŊTD���ol��4L<v���[\��E��=�W�f���!j��3�M�8��2��b�g7P��0vȓs���i��Yq�G�֒�u��]�J�rκ������ؿ�L�&�m�>{3v�r�6[h��1��`:��n6�Zo`�#.-P�d^���<��sx�ߋ�.��j�j���&�����%�����0��ce��ng�ֲ���Դ�y[����^j���Vo�2�2��evΒ�T-z�ǐƾ�;��- �<�WO��sg�E�[�{�ڻ�RѰ4k�D�lr�����'�i,�u}s;��ۻ��*�Q`��q���g��"�@���޵,����ت�ֳ���!V�ERJ�٥��A"<�m�qo�U4[d_ˁ��
tē�e.�X?���C�x�Ymg��;nяt�����K�Xn�T e���e��Ϟ9���M�ٷ,h��Mf�A[��"?Á������h�����|��2� ���WJE��)�W��Y�� �#2+l>��vXV�[��&]*>ӫ �H4���y�W���?l��-���{fI)\��	9%L���_FIV�R�N�I�<��}q"�Vr��Z�t,j��T�7�B�֙�9p�)C#Z����lp�Z�#��`�-=��{�l,���Ң��9�M��/�J:X@N�T~~��������\���T���Y�
�{#36����.�a&tÈ��Y�#�&��E��8g��o�I3~o{C��v������ê=PB�f��� u�l�K
܃�����Q��{V[���୸��r�I.�ogg��{���t�,��a��o�^�c��DX�pi���e��;3�xai�L�y�D�C�"���S.�~�O�m,6˸��2n��?S���vF?�/���ck����W�ѿ|MC1��E��ELsU���I�����֠t�~kޘv1�L�d�K�^@{���YT���{x/
�K��A\1��r�r��v8}�&�Iq�p��c¢�1�?�U�M16�� �0��g�\���%,-Z�U��U�4�>x㙵W�U�C��摤�h��
o.�7	�'S���    IDATʲs�Ņg.`����-�X�� �]k�|}�Gxǰ�
�9\8{�/_�fwW�[��{���G�������6uX��&|?�UW����,:��S�w�����C�J��]���M��]H�*4\,xGfLQ��@&�����"����?^��f�W�����S6mrB9L�R�Ow�j�CfA��<e%DF��N5y��E��E����Jj������WK���F1���=e���Y)ı��MM�#�%�Av
a�Dr�3�TN��&��@O��w#z�����$U$���Hi��w�Y�y�?��];9	��!׻RASן-.^�X��-��PB�.�^ @΃�܌����].7��3g���݋���j^t׍�ȧ��ϔ�C��t�}��1e�I�}h��������{�+��Ϟ9+�vw�f5�Qw���DX�����p<��}��a���?���h���>C�f�	ī��9����}���i�mo{�^{�%�n>���G6~>��'p��~a��ă8��6����������Mi��n~�ϋ�\�2cȣ{��s�ٗ,-/�ߕ�=(7��W�h�
���)�&�ve��bB��M��U�,�:��R]ۥ�t-����j6{x�i{��� V�Ec�ԫ٬���PL�B����X 3f�I<[Z.�'Uv.����z�<u
��V�J�b{���R��ު��kζj�<j�#O���q���wqic=aVT�u��uw�kw۪��휩7>��b�8w��~�����Q�|�F�ZM����.=�1A+k6��{�#AqҪ�2�L1ۯ��as���cm��{a�����!o��8+L�4k�-<;���3}f�r�e3�5��C,7�l,�?�ء\���YZ���ƛ��v �u㊍~��:��D�ҋqq�L&'MI;����M����ct����,�Ǡ��f�A�g����;�[2 ��'��T���sk����E���ZձH����.U!�;
�ܼm?ݐq,ؘ<�k�£��1ն���T��}��>�?�����꿿�ն#��w���:���������v��Xl��n�k��R�>��w��wP���Pp4`m}C�$!��4��ם`��ꙥ�,�Kxꙋ��}�n(5�&����3ԗj*f�(�hT}�<,��_{#�ك�7��5µ:��g8�T��B�cx�廳�;�U
�ا���=#cx{T�p:��A&�U��e����#F@w�#ŭ��6�ٿO�H��/h���P�Վ�1h��Ae�1:�],�,	?f�V�RT��`o��j�e]u�N^رl$�n$�#J �0lu�P��,S�I�I�pr	��SF�ڗ�Y�6Q���z�yy��6QmT� i,�����ٷ���%4EZ]רG���ߞ9{G�����q�U��?�	��c��<���Ku��� ��{Ntȧ�|R��y=��:(��SB$,Ƅ3�Fo/<���qkʲ�3���;�7��FK
G�՟�xܤ_rb��b6o.O�Z���l��Rj�,�s)��4M��|G`M�v��\{uޜ|�l�j|P�$1U�{��jY�<\ BS��T�$2��x#�Pw�f��R�K�'�~�¬�1ρ"�m�X6k���y�]���5���	���DE)��q�pq�����T�#��ډ$�dlqL0nO&T+�ą)��[�d���]YG����+eS�H7�`k��N�������~���]o{=^u�q,��|i/�}k�����'��������m<��%2{�D�����s��������%'p�PtFK��/]��D	�U�M5��!����vq��!DF�!>������i�'y�k�tr�(G}�}�����>A�6��}˸󎓸��>�xC���ٸC�t��z�4�c����Fq��6ݐr����l��j������H�K����Ϳ5�l��lZ}rl4����N��(Ǌ�X�d�6�+�la��t(�1C)T����v�)�Y a8a�ohg��^P��/+!z#�cUk�{ee�P���PԘjŷ���֤u�@9�o��G����n�
LU��bC���\��T�յ�A��=���Þtȏ�8��V�\�xQ�5��89�(p���������u�����7��m=6P�st�C��S���r{��,�����g�_�n�}_��8��#i���Z����A�g*@6N�/�l����s���;B���tQ������PI�fk4��"&�_�(w�X�N�+�2�e�w��D�"�,8��,��(xk,�K���}�32�����V��i(Rta��\ո�v_��<p��辣��PD�>ThW&��52���s��i�b�����dx��<�"��$	 9D�&Ɵ�s}��t���'O��O��[�����믑������8t�����S������7
�q��S�*��/��%c^���~��kO�.�_��mҗ�O�p�:�?ZQ?e'"�a�R����)u����!���g��*�L�o^$�K]63�a`���xΞ[��7�E��:�x#����RJ��}<��p��)�O��cY��>� ��SO������/>��~��%,��#w�s^���-�E�5�Gh�|�Q��$�\�gV�� �|�)�y���ءZƩAKv�%� ���4l,�a���|�`�%E;�h��hWf��W�:�U��[W#��)euoᕔ�Q����\5y
≢�)��m�����O�!)G�[���>q'�m�\AUB*(��Е�V��xMl~{{KA{0�0kcH��[��.�]��3���[n���
*�&Պ�)�B*�1ڶ�Q�N�7n���̸��L�+�f��U��1ī���ɯ��=Y�x,T���(`���r��gӦ��?���;�g�;�o�Lں�����#��GMÂ�QsG��fH���ٌ�zb?�d��B�����]����~�"�p��	�X�?%\>�6l8���d��"Z]n�J��P	g}ς���`Aʳ��X���cO���2���0T����hˑ�M�#�4�3$�sR���!F�6j�3�������S����k:w~�,��"G;v >p���Xl�|�R�Z�"a���=���}�瞻l+9����E�B���6|4(`/��7��Ձ��,�\�X���O?�g�����/`}s*+2Cb̳>re֥�x��o�/�-xͫN�� �(W���jSt�v���]��&� ���?�׼�N�GS��>�3�;�X����=w�7��|��+c�Q��������=���:&��
�0Ȏ��[+�����:W�1o�#�,}Fqn��[˔Ť��HO��5�T+�H����YK�:U��F;n��^3Q�(��vǄg�hC��B^�	�K`�L���r]������6R�M�R��G�����2���s�tٶ�̲m��6R^o�>�y:����L] ��k}j�xSQ�Gb��#��?�L�*z��ӈMC��gɦ�t[͙��H��"_�]6�R�d��v�0��Y��w�~��<�<3�TWϸ������lp�W��h�������� �TFVE��eAe���4&�es)�Ŀ�|�k	m͜��8��\�Yd7�o�Y��g�{��j�>.o�;��qRk�0ﲭ:�u{st#h�F�w\�|%�w;��o�eAZ��K#�sG.ȶ�_ب�c�s��)B��n�{�E���o�����>)����8��9��U/�ٳ������#<�����������hE��4��M�t`��7^���u3N�ڃ���u��_ln�8��D�LR�ݳ�"q*����:�?������;��˛���d�Ҽ�a��r��B�����~�m��W� I ��C{Xi��M*���6�s<ڐr��D���-!����O��o��z�0��������ʴ�S �5�-\�:Ύ������2��,����>�G�AI��������4)���v����7�BW�F手���"k��E�Z�F�ӗ��[��=��m�Z�J^�����z��yVπ]��QoU�Ǥ׶w�2���7�`X�fe~\3���&�JGl+�F}ɦ�	i��-��ҩ�l��d��r�����*H7������󷓢��c0|5ntif��6}ծ�H봾�X��`M��D斋P
��� �:�H��.�2�؇
rk"�a�3��\�;�����X��u���F*�2��hPu$��75��hV�,Z��a�\V�!�M���9[0�Z�C�EX/�Xw!���<u�0�`̊�����-��,^���w�\���dN�?鑊�QDKP.;�`W�
��3}|Fd�ٵ=�9�#�}�ƼT�s����v���v���y����'�����S����/�������-���g�?�-�z��3s|���������0�t�\�c��"^t�5x���ͻު�En�������&�$��	�=�h5�z��<~�=�_|V��3���ob0��FJ``CZ'�񶯥�����WތE�铽�� �����'l�+��n{{���ؿ?z��FB=�y,>D>��!��k����~��a4JK������7�lX82۷�n�kٶ2)nU}��MoD���V��D�^���mX�v�d�|6#�Z�HB��LP�����^)3�{�K�T��ܾ`�	74iYn��D$'�m��p��-}�JlW��U�i��	>G���;�2�"
������q+Z&4D��a_��ڰq��k���+r�T �̖���X����⼀����s���9[XK����'8� TdU��L��,��Ҍ/�������*k1f�.m�^DB^vZ��a3f?bg\�,�vu��F gW�v��g<OI�6�^[���lJ���*ϝ�cH�I��;o}sw����fbm��Y�_����/]�iE%(�j�,��z �& �9����=}����\�����,f�=/�}D� U_L9���z�:!vKg�J��N�"�c9�'�|&9�:=�w6q�-��]��z��a�
�������~���.��?����9����;��~���������zss�i�.�����w�t��UcM{���7�F��?[��LV,K�Qk�V#�h/{�����
�>y^�p�Yc��Ί
c2���r����D`�^ex��HA�UȒIV�r8w��t:�r8~�8�x�	9rDcbuu��-�Ci��8���w���øOZ�A�n{�{�f��<�Ja�]���0��Ev�k��ov�&E��9dv��ae�h>@�K�JZ���`6��u�ٯm>+�3����,�yN����M��Ҽ��
O.8�j;v2�p��FHE�TǓ#�=ev=���X�Ԕ%��Gܘ��;k�Rd���-,�mr�7/l
��mk�%�bM��N>`5Bp��S�p�J�My��Y�����(��7\pC�+x�~J^)Ğ� iw7�
�n5ѸM����M$�p�q�a2�?��J�o2`C�� �Q#0Zq��l�Nq�T
�rDJ���N�`H�ߤ�I��N��SC��h4=��;%f���H��m�#ѧIR(�}B|"����c��$�L9v��@P�|��{�Ə�A@��CE��=V[�����.�1���g��$���)u$�mB06�Jի"��g{O��	ڙ����7���O?�} Z��~�q��*:[�~��� ?�S?�G{�}�7������^�����v�{���r��8b��b��Ag��tXMw��ߑ>Nf�E�ލ���e�|76�XZn���B4�c�>��=tF�j{�:��Xt1��et��d�����dLc����9䦢6�G�䝝��]zu���`0�\&�x��\C���y�巽�7�
���A1WC������%T$P#�A�D�@1.�H\�
�j����a�!�K��9Κ`|��W.�^53l���6ւ��`*@z']Zه��E���AA&�nQ�&� ���9���5|PJhF�A���F�c�
�95)��W4�k. \����*>䐩�4bQ��th�	7a�\�@�Y��j��C�Q����mg�;qMvC~p�}b�X��lP��Թ1���ћ��`�b�Ad:��5:��L2��WW�J_���-�W�`��r,]�U�a�����2���g�pT&�����P.�ϖ�{&랔aq��Ffm���S&��J�A_����bh��;G�<;?/�zW��B�8������u/�f���IYK���I�fL4Lg��5�%J#�� eE�^FA�Ϸ$&O�,
^�=Wc����ŎZ�9�����e@�����4kM�m�\�L.r���f����Zn���V)�ԩU����D<��G�;n�����<��9\Z[ǫ�~�ͱ�_����}�G�;A�^��bCދb�L�����p��7�mo�F;��Ol�ԩ�͙ �|�\�}�x��ÿ�����~���я�~������Q�攈a�v�[ؿ4�^���շc�bQ�|^yB��L/^��~��V�%��m�1����.���7�l�6�L,�4ZY?�����.�=�u���M�0����ܲXހ�?<bC�J�~dR`b6�#�&����l0��\�Y��9��.
$̗�԰.e���0��� �E���|���>�C��Ё�(��n����Ŋ̌�l'���/&��O\*�8������~i]'A[��=Z�]^��1vwwL6�v@�f�G2h3�}��.buϊ��7n����ټe��6��-<{�y���������٨���g�8���b������}٧ydZ�EG�ȶ�i��`���V+�`�����gfs�$G|��=4� >k�w?Rm�E�kh�V4�|�D��z���B8.��G?��9�AQ�}��\Y�
��i'��D�rμ��H*��i�m�	���1�˶�7W��4���=%<4���w'����2��i����/8�`lψv\S�"�xQ@�?q��3$An#a������l�7�NՇ�t~���n�Q:�M|�7�P?��~=.�m"7���UI���8I�������y|��_��	E����p6�'m�fY��7�0po�����z�8������8�.�����̅.�<������$*-���A��<�Q��B��Y�����N��'�4��?�6�v�bE� U�df����� qXi�?2mf�K��L�s/,,��a��E�� ��Y���}�p�BՂv#�����1�H�.O34IB��[�Y8�g6���
�VB�|�����VLX�ߛ&�D����M�@�*,i��;&���y<�Y�-a���z�e�t��¦���Fe�Ov�l?�슎���8�!��0{��tQg�� l�#\�1�����G�y���7y�;���u��� �Ͱ�������jbq���=�&������fϗ�&1�RRmn�^¹3�am{�Ğ}�q�mw��o��7((���.�N���~����-H�*56����m�ڧg�~�`�n�&�;Xp��o�2��6�DfJ؄�5�ħd�Vc�@fku~��}�&��Y�(���HZ�1EJ��Kg y�_��=[��w,V��?���x#�L�@W=��bcL�<W��(�
��l������������>'���}�Q����3���m�>�Mr�YV��PEU��XE�������˲"���yL�l���t�������7vq�icl|�C����O��L�Z(���G�ݸtqk��8z�Fl������-G�d2�p��
�)�P��ݱ�x��ݎ'.m���O�{��i��/�w>y���%�ˆs,.]�B��q���%426����|��q�uqñj��ԍ�6Y2�FX��H(�L\�c���Cs�PP��w/.*���.��ϟ����{�����:rw��}sRT�a�{C춷Q���Zlb}�"���F@����C#.w!�^R����G�b���lb�|m��������k�,u�g���e��>���3������G��rC��Y�(S�1+�b��X��\d�%�X�v�$ćI �rn�@Z��s��<��7\/�nee�z�&5N,Tml� @࿡��#���F�`���mL�    IDAT�`7�6�p��<x��o:̴��v^B4�D�T��Sc0�'A{��[.�n�y�J5\^�T���LVv�O1��}���
O�z��
ݟ��o6h[B�B�$,:�l}�%U�p�X�t�q.,w*���z���EHw�I����/��v�<�HS�[�c]��df���wcXA��D��Z�	�>�;��X��P0t������	F�2�w��^��A;�����C��?�`���2$`3p__�g�9ǵ�P��Wz3�)��x{>v"���l�����t��6j�%
gU�I�3���K&������o��/=�/|�s8u�Q|�����5��?�8~�ޅ������{�M�����4W�Q�c<J��D�Z�I�4�G3T��P��6c4�TW�8�SAexG�=��/�Q�1OP_9�b��b8�v�P$2��C������ux�'����u�O�����)Q6���� ����1���V�ٵ��f��޽��+�r����/��_����g6�{�[����{���b"���q���)�9~\��+ut��84�20��#�Bg�
�dL�3���xd�LIac�b�Hj��`��Y���9sX9r�����%X�.��X#��mu�Դ@њ��\E�	�:�0F��M�+
_G��,����<��e���XG�VG{w�ј�vV�x�4[L`�㭧n�<+�{b�|�&���Y��)���'���6��N��6����8r�
<������S�2_-)pk �ue�J�h�9lt�+LC�y�����5 ϲ-@�]�+?'�%OR@���P��x*�L�%�E���1�`��&D���������d�~}8�S"	�jxI�j��̡�$X³Yǫ5^8$��b��L��K��]�CQ�u슸h3h+�;+��ĂL|�O-2���|�N����\�����%����/�*�U�L\�d�F�)w��5��s�nM:���]�kIV�ߒP�v����M���v���_�^{��&��۾gO?�0�xً��?�n������c�w?�_���_�c��
�����^{�%f-LGC�TGj�3�#��->�{��i�0�Sn�2b�MG�
�+��`��{N�U�����㮗ފ{^�2�����y`�M�2̀�u[��Bs�t�;�c�&��7(�e�#��U�>��$����y�}�l�Bn���˸t��0��N�����K˸��;Pk4��v{,�Y�i�ZWT��n�*���i@��!OL�ŋ��^bA�eS�96]�����Z��去T�;r�Z�rL9�,�"�uM1�:��eb1��<*���H��
#��vq��._���O�t������B��*4��NW�˝6�mb��oi����~��G����a]^�p���A4�mP67���lm����j%>rͅ����j-���s���X�2*��(7�2d�����;�t?�������#yu�u8�.����;n��NS�m�iN��"�X���{0��m��d(��Xۅ��������e�p��-[\u�e��-+�Ͳ!2��b�Iӭ~`sP��'q����"bd��ff�ʴ���e�)�$b�i�3�P��B�12�L}B���~y*|��-I���+(�6<���/�tyw�w.��E��n��H�A
LG&0�l�4����˫�י ]�IU���[�=�(7�����G��������k��z��C�#�a���j�'#r�Ji	��1��.���;�I햙���b��A$���&J�z�'�.#7��"�K�������lz��tBM����E��T̢�4���8a�ŸI�={�+`s�����8N����C��=�zr�x�oXbѵ���?�qw7��� �n�	�+{�q��ɔY�M��'p_�2L�}�߭,�ۮ��m�t�>�8�,�g�aт�����Q0��;XZha���%+T����>1�Y�6�� e�r�f��ϱ��A�X�p�m������Ǝ�{V�UD��d���RKm�\j�v;�i�Tt�~0k������X^]B�8���"��m���H���M�yT
�k%z}��l������A_��_'�jj�y���>ϡ�㖍���� ң@;����U@O��<�
* S��@��&����SC��V�`��Mv�'�\�]U LÖb[�a�mE�̅�)]�S��se�d���߆�[��Gb��P�lƝA�Gʗ'��E�.����Vʌ���U0E�_{��݄�=�K�.�8w�%��Q;���u�rwB�i���5-(���-��l�C&3L��8��\y�"���7j2�pQL;1��P̊�v7�f9l{�=o-�~�M���c�d���M�ܳ_��NY�mtl>nv1�5��?�Zs��j�z�us$����0��Xi�m���E.��XF�Sk�]�|������61��f��. ���g}�ؓ��'o����Ts�� Y�UlW��]�'ZA�嘏��}� ���B�P��O����A��G.`�/ w�7���T����{K�&���Z��]{�+�XZ1ݍ\���L&W��@el3�Ƅ1"�k�7/5V�MӁ��l;���$�jU�풝a����T�T��']�m7.3
є
T�� ,c�(�G�`s���w��N7d�t���k����贻���ᱴ����\�r0;�fEln�EK��55�]m�Z������Rk;3t͡<g�I`�3��5\�|ǎñk��ڨ)`4�d��h�f��uBS%�175IS��	��lS��O���Z���z��0M�?g�$�[vݕ�>�S٥W��Y�Ċ��}�`�W�op�=�eM���Y�T\_�x3Z)����	4ޮ
�ᶓ��Y��ӹ(I�{�;��L�Kx�Y����`2e1�G�o����N,v'�ifL)Zvs��nF�@��Kتe*���ž�2hǂ��f�ΰ�x��\�M�H�c��!����f��HW���d4E��Ǩ����%���]�].�c�U�C~V���7�Q�Q��AX�O ��/�܇B�;�4���H0�(^��=d��h�ʒ��>��4�e��Xn�1��\�s��z���d 1�( ��.b0�軈��9,�
��e��_�9PA��=�*x�������4i��*���-
<������d^I\�D�.�M���s<��:���Ƚ���W3ѬK�)�y�i} ����b0�P��D��J�a��Y����"j=&#YD��vtʡ��/U�fv@�����O�D[ ֙5),4[�zG�`�����m�|���ϋ��u}Ȁc�|h̬WW��=���Z�A�TSk����q26}m鎐�r��~f�U>P��KET�#+�
?#��'�m�ѵE+����άY)��6_I=0n$HTg�����E�˳�V����� �i.��1�;Ȯ��KY����ht5'9�����-�k��&�v)c%�Rf\�d��BQ�L#nCK��!w|����H�f�|O�e>ԖV3��@�<��eS�vi}$K�K��n����z*�p��#>�,8WH2�����A;�E��l�kTz�j}�|p�8���g�p��=9��xSL0\� ��J��%^���B����d��P��v�l~V�t�aN�3��Ř����#i���OnT�?���ùӗ�ll��_cz�'o��_���E<���^���y�OKoga��&*�*j�:BF��V9O;��60��P���}��Ml)c�B���m7�S����墤�5�fCA0�	M|ٯA笾�[��6
���ƻq׋o��?`nP>�W��H������X`$D����v�����X� ����;�?��ݿ�Ǹxa�������,�4U{=���ml�\©�nW�5}�h<�+��!����7���G=�3������9���R�$��>;��>8�	����=+­HţA&���m�/!o��-�zg���&GЖ��h\jkW��N��X5��3���h-/f����;�!��U��z��zD戏��l���p�`��7'c�����U�
�����'Q%F�fO��
���>L�wg=۠���Q"��z����֓&�Db��������E��,�M������L�=�ɂ�������{m���b�dI $e��.=�C�ӿst�آ��ڥ](*-�Y�(xjIO�r�d�yк�ƦݎGo�'v��T<e��^F��gM��$�מ�Z`�F��5Y����I�MIE2����1�NP�Ғrf�/Ȓh����0�H"��~�V
0�*j )�E���#/,��o�ި]$�Ntp�YV��"��&���u��8�W�z���p�Q�|�~���DW�7��?·���x�gp��[��C%ܴձ9��Y
6����ZM��4�f�h��df-Z��;����G��������n��<�L�^sg���y�>�˘�}�	�
5�7)���ģQ���Jw�v�y���ݨ=�x�;;m=��p���ב�ϚZ�>���n���J��ѫY���V�a�����~
�������U�:��8|h���sg��琬uFj��	1����VN���%3аuٚO"�#l`�Oƒ�>��/�t�l;��?[I�V���d3f7�����-!5�(�CA%�
i%���#]f��#Zu4t}v��������Ԋ���@�5�(4�9̥�G���آ�g0&��N������vاP�)T�*�P��_A�ҚN��f�`�ZB�L���q���dPiqb�>�^��f��)!��:�%�O*�!�t�v=���?�o"+�� �==�V&�aAH����h��f��x?�]�-��5�g�=���N@MBl0��I@6#�¦�s��!'}�WfԔԽ:`_�OG�TǦ�4�%��
+�M<[qe'9ϟ:+��{!l�-2��k�8�����u`���%
qH�A�y/+�Jw �<�N:'=�kHwov}�_������i$5<������:�i���?��o��>�Y�ؿ�V-����G���3��Xp~��Y�F��e�`8��c7)H��i����f�c:��_�����.�u�xN��ġ}%9��J~�^p�A|������E���c�N@����&&5g�������kW�i_��t����zk�v���M��p۰|.a��k;��>�-��N�H��ϟ�@�4��?� �|zhA�i�jU5���,���j%�1�n��ɢW
��ea`�`b�
�p��S4�o��+��U�
��lٵS/���v��~~v#��R��Ly�'܆�U�\�xdE,bJ�31%7��){���ٌ�d�P��ʭ�
�=TI�f�N��rղ5�Lfr�׀��g����P�*�\�cMdI����)�nf�����=V����&42�69�P�)�H�Ԋ����&ۢ�`�'�"���W��l���6G��"�d��ī2Z��/XWg��@}�葒Q��u;fdP�r$��D)YB�}�F��l��(2+Fz�Wq��j��:��*[�TB�Kߦ%�����b���,K��].p��hm�|�ݟ�.4�<;g���Կ����盵G��'vU��y�����a�+�p��:(���ݮ̴�;b��O�OS�7�|>_�0W89Q�zg{K�)�����7����M��>�������ƥ1�x�9\s�z��U_�~��x�ً���7�ba����D��α������^cY2���߃e֑op�'�#_��7Ο>��/�o���|��ǭX^;�)��@ƜA {U��kN�ؑ^r����M��jl���1O���;5�x�⺑(��'W4�zk�*�<IQ���q�no����ছ���/٢�{p����9�t�C]>�UU[�7QKk��5��Q�͝��y�,�z��s��4�T���4#*`q�M=ޜ"'����ǥ"l�8Ū�
�\q�QV.�SH�^�RoV1����Jm��$�o����w��M�d5{��=�Iĸ�ư���pq��+��εZ�!7�a4�>���ǜ2]LgeL�\7�!_���MI��N�/�P����Mv��	'#����r��eE��|�^F
��c�y�(�e�;�j%l�4SJ�F3�{0����{�- �#�� #��x�^��c�4�0��E$&���h%L�Y}��s�E�bq��1�Ɠ��f��d_��m`��}��}��mY���e��Ľ&���xo����}��fNj�[��p�X5��:��Ů��᝔Z���m�Pw�v�W��v{L����(��htd����?��;R��*$�|�J;kg��v	�/���Z|�^��St�s����c7����7�V�����7�'O���]��$(���%Y��.��-/��?� �߇o��5��xu[MuM��A%^س�B����
ub����ş{����G��J������Q-�p�5Ʒ��<��'�o�F��SR�	66Ƣ����R���R�40v�T��ٵ�D�Vr��TP�gQ`R�c�?��cm����1�W�{�׽�\{�3��Y�q�f?��c�=O�1����ڰVU��d�]�sE��h;����@�ϰC���p�fEv��I���8��,rE-Ps�o2��2�[��!*�U�4	7� �5���Kd>�Mx^f���f$D�36�bH݃"5X�S�*f�1�\�g�W�*`�i6A�g�t0&RT�7��G��:����c:a��Рa|��E��x��}{T#`�f���4�Ի�v���ϊ�-����m�6K�	�Q��N�+�O���i�0�M����p�6�Q�K%͚�,�A�;�"c|�����pn_P���2@%������j�W�������H���W�Z�����UYv6`k�g=S�݇�� �X]f5��a�Y �%V ԥNUf�%/����h�����k"���{�ǅ�=�����x�n�+��)���BAC􌚻�`O�2�k삖Y���j)��̈�@�4F�%G�h�ݽ��=oƟ�{~��ߩE^�t�L�|�������7\�<���9�g����;/��X0Q�<a�.n�~vw������{'���(�%`�.�*�/_ƼX���e\:/z�KQi���
_`��9��_�]T*-��d� S֎�}��Z����N��=t����۵Hq��\,�P�����܀�Ta����ݢ�ƆҒCgcJ��}L�����̓��ӏ�|��U�Z`���y!7���u�h�ֈ�v-mؘ0�Ur����4*�	�p5���ݘG�;��0�X���`���G.��'�Sq�j�aC�ZY��A�Ke0f�9�����Rn�F���li���h`]t,tF꣦���@6g�0JR��l����3��1�� �c4e�����%�pbٴ@b�.Q�<H�玂��Bm�г��P����r����Asq��i8b]��u~��K�C��fp�5Y�ט1�(\��;ڒ�,�U�u�� /��i�t�� ���b0Nt������sD��Z�3��� \�_El��)v����s�@|��F߾���1���*,��̛����ų�b��X~�gR )�9D��l��U'İ�o�l�>��/��lT��W���+���S:��"���g�'��~.�
����f�Oubǌ���?3�C0�)�d<�W���|��n�"����L�>�������&�����?�Nl\^��, r�����Js�rg�<�O|�~��k���˿���|�s2讖)&���S7^��{��*<��ť<*3��(�x�/(�:v�z<���+�Q_����w��`4�q���?�����=��buY]���s�DnԋXZjH~�moyN_T�Ν	���
��la�A�`�Hd��1�tj�El���[������h�j��_�}�Sf<W���W��{�7��|>����oR܈�r|�j�fm�cK���j�
rT䖴�-��[��ܪ�;��¥�>��N�=�2��7�����;;��pef�6~7כ�Ô'��� �N�[�h�ϒ{Ɂϕ����\Ir/     IDAT�ފoi�u��ٞ[�*���@�aN�	oş��W�T���Fh5���p��E}���9��v��5E��Vq��6�C㰏�P�V���Ҽ�a�8V��m�,�='����Yoo�v���"3�B���6l^%'�s�yI&�Ik�OzP6M�i�e���bo��l4�x���Z�|7#xLTt�ad����5��N�e?5��.�5��_3{�@f�XE�V�ݾ�ܔ-f�'X!��h�g:Cy?R<��g`��t�<���!d�������az�|�v�|��C�����\_]^����,r�����-"U����O�I�u̲w���	�I���C1�baV��NNt�4s��Cg{��6~��>f�.>����[O�O����_���g��~f?�}���_��c��[x��M�Īe�ؘP+Z�����}�e���z�Ϋ���᾽�dD �f�;�>�����IT��ú���?������0n�?����W;�I�����6n<qH&-o|ëq�u��"�b�!�������Bj�5��f�ϫ�)r�r���]\<��#_~��YL���+@Azگ�5Y;3hת�X,!����uD���k���� �b����]�%9#�Y&U���<�@zd��/o��gL%kyي�>{����~�;�
^�L�Q�k����m�.2�*��)���1D�ɩ�+:��iך��#(k�(�����ԙ�0-�8!
T쌚�V$�4�-7���N]��ڷ�Ņ*.^����7���M����b�.Z��ϵѬ�Q�r�L�=�c�B�6)Y�f;�G�ۛ��X�pեe<w�,�9rן<i��j1��m��F N���f]l�A��Z�Dd4ed�V��������en����jr���Y�>[�?k�N|3�S~���!A�
�-(sR��Z����
�?*�{P�kA�0��I\�c�(,'�ϳ`h|��P�M�g[ğ2jv)vW�F(V&�����g��.mky���l@X�/�
� �q���+�ř��,�D�ԟ��a�y��d�5[���ƀF�p�H���p��[�Zh��6�ix�F�	ڗ�n=����K�t�(��������u�ջ�?�_�;�����N����طrJ��c�]��5�6iT� M1����ǫ_u^���Z(�Rd�h�������n{��ܹ�%�Z�װ������XZ\B�nP	���>�9\8��|�v������y��8:c�|��/����W�#-�=����U���܃�^�@�W��$�bLOX�U�;C<��G��O?�/>�Ɯ
�|k��Yو	��A�^|�o�K��E�1ګ}nŊE��|D��<��1�b-�j���v1�;^�/=��Z���'��#�r���>�o��n���]�b8}քU�K5<��.l��=�<��a0��� �D9V�)"4G�4Gwf��UB4��Z�?�5��6Q��.�R���3�!��)�.�0� 3/�^-����Ѫ�P��h���G[���8vxvߣ�;8̅j�����)�����؛@I�]U��������3"32rϬ���Ҋ�JkkA% �hZꦛ�A��{�{�=�6�g�A�,�
��B%�TU�Z2+�r_b��=|777�����gJ�c:G�-����}��+�e{~9_��VG�ލ&�C؊Oe��������U�;w٪RK�<n��viZ�l���k �4����y���Bs��f�MPc�ٛ�(-�/����E-6��[��	M��I+*p���D�׈$�(\�Y'�g؅��2=W�^
m�~	*B�c6��M��|5��f��m�������k��0-�<R����#�t��,^_b)��PHN�r�UN���%�m�4?�&�6���֌�m�c
+Ui���@%#�����:��bCT�X���H�|���X�|ɶ��:�h���EkgQ�F1�`��%Ѣ~����7�7�/��������U��b�ů��'�O?���o
_}�%$Q�ɹI9J*o�{���G�1���9�v��R���ƗL��a)���"�:�� ���,�P��P*�͖p��
����8y�9,���u�H��Gw�uI��4�mn�;UL����o{D~n6[8�oR����aI���psRl�7;X\��w~���\�x����df����/�a|��p����O;TR�
6)h���|�!��d��͞H/>p�f���>�C�>��E��]������� M��\d����fHG��.m�}��Vqe����x��Ǌ��."4��̪E�����*�C���L[�i�m�\����(ޭ[2^F���D�����ڥ`�w��v����w%h�	�L ���
�r���ն��ͭl7�x��JA�*�siy�>6��;Z�_����^~�6��"W(��m~����
%t�M�*%�Vb��u8�b�����=1O7y(�A~Ji{ޣf��+k��hx����"�|��gep�A���ŗ��[��@6���&2�s�'h�lV/�J���X�h�3eb�?�e��a�Tz/��ߌ����ѐ���Z)�����T��TD��ٵ]Dl��D�, �X�͍7��+�#����T�g�g�i�gdtWD��,�zmT��ل�Fw�������g�
�d�PȌ�4�$6~�V#LON�7�tܚqeY.֍�=h�W����y|��~�m����Y�������-S}���^Y�x�`���?�����ULMOcWe���������>$m��#rvp}qQ�p<r��`�1�^	:��ٽ��!sc��?�o�i<\kWč���ESK����Q*w�{��\:��'��Dn�P��� �UmJe�|��%�4"\[��ן:���C�-"�%�}��]�^~���m�\S$/�y��ҏv�1Ӱ�L����®=J߻7���v�+�k8�w��`g��8\��m����@��6�	�خk@�����-����F�@#�Y�v�i�j^�T�R���T&��p�l�a��v#I�6����	%��|쪔a��'�Z]�I}|����7=|"��D��$P�a7BP�1;UA�¢D�K�tu	����M$���Z�"f*Y�����]J�F��n�n�G}cĳ�~�	�����bbJ�m��\zl�.�1'��.�*�Cn3ŭ�	��n{X��9���Q����$Q��o�,SU��4k$[�`�t��/�;�)
~m`{~R��?�oⰲ���5�5A �84r���r���o�@E�Cj���A�����U��x�⽄���jq�!at7g�u�J��s���U��A��ֺY�-S�Sh�%�f��D�F�7�ċ��ɶ�2��	m�ՀV�>g�&B���Q�H�	�/E��i�B8E#_�z�w[�5T�o᡻o�{��y���O��_����������)������������q��A�=��Z?񓿆ru�*AB��O�g?�~���EC�/��I��F�Ks�s'G��GvX�TB�XD�+�׉��?�,���:��G�6��"��Bu��n�V�t.��9쪖q��.	�ĶO�<�}���zg�ښR�.]Y������x��� �8�^��\�<l�!���JiJj�Ox�{�\��qh�AQj���r|Bv���9�ޅ�܇ބZ����"N�?�[��	�4v��w��o�!k��lA�>��N���6./�x=t�6vؤ#]���W�����0�&��t�$\G/6�e՜�c ��m��ݔ4��/��}U��k���Y�A�����uq��b���#s���x9Z5P�\E&��ǝ�5���Tߛ��v�fsO~�$6�k��ȏ�߉S�7�ؿg����PW*�%ȗ�$hwZ],_�����hl]��M��(U*��G��Fif2mÒ`͠1�c�!�Z��*k�pS��A0�,L*A���� ���d�Z�X�!��\�i/��lQ�i����DV�D>3�MTa+sce���`��-H��H:�o��d�V���I�K�IT8I�����kQ�)R*�>s�����:2RHe�``^����Q�Z�Gm�,���\a�#���HMV鞊�(�I�#h�=onZe� ����0��c�;#���Ѵ#�G�a���/}!��V���	��ƿp�������w헬������>�Z����ceU3�������Џavw�/v��O?����K��c�p^��� G������xE�w�;��"�Kʤ.\�x�X�Ν�{�fk�˧�au�����/��ˉ�_�Oݗ<�)$����$����ݎ@0<^q�^Q}�Cw����wWW��]?���9�{�<�����O�C�G3`���� [P�1q�D�D�Jin q�p�}��%93S�nN,��~ ]0B��H��!��0�k�>|¨������6�f3���a���/~K��:5�(�Ae|fv�E&�G���|u�+���l������>��:D�ti�N4y`�z�R�8�"�F��r�
�I�I��`C�z-��BL3	�ʆ(y�m�B�K�kr�;�؇�G5���]D]Y d��kW��v��ơ�n��wE�0�i��ٗ�ſ�*<��خy���'Ǒ/��ޒ��dq� /���Ύ,j[���,��(��hd�h�ͱ:�?L�kd2�ji˽�!����+R3Q]�Y�.8��� �� �����u�>�}*�)]x$���-��|�8�h��8�dx&&K�gZ�������P�8��������q�cU��a8׶�X�;UT��d���7��a})�)XN���t?�L(�%��uuj�ӛ�-��`����C)��c;�a�2kb�@6�Q6��9������7��
�𰉏�nY2Bk2~O��\�@(�l]t��;���}e79�.^������?�><����}����}�z������~��x��3h4��_�)�]�����J�F�u��~X�K�B��g��k��j�޴?���MQm4����������-�xnA���F�W���^ß~��بsG�2Y$\ܸS�sưE�L(�@Ѝ&�R��ѽ����ɱ,��F����W��zׯob��CK�d����˳���(�E+���T�G)?	RTe:�����9�ą�x�.Z^�F��G�~���s�{����x��}+%H�[�I�w�����M9���O�B���$~��;�b^^9��_P������2~E0���Џ��7��ק䠈�g�q��3��L��n�����[��4 xf� �mÞm�ww�>��É�3p���nnb��U�����t"����C�����3��Eqx���>�^�v��3�ڥ֕m�l`��6��5��ctJ���Yk���y�v%�&�͙�wT1d 4Q1ŋo���{Lvh]U��i���g����Lmʘ��5e1�y�1"��h!͸���n�0u��̬6?Y�eǘ�4#��	��y���7�4��Y���
�g2q�B�.�u�\M������j& �)�dS7�S�d��H����.JN*�n͚D���B(0�֌t*��'�Lf�9���Y_��'��r��=\�Y8%sH��B�M���?t62��CR�j�U�H҆y�d�9	��;�4Np��E�֯�+T� ǎ/�]�Ns�����|�k�09Uű���}�����gq�"��?�^>�'���i�5:�|O��1������Ms���D���hL(،'� Q�sǉQ-���\�����~��?.T@�A�(+���>w�.r���&�=FQ�"�!4�$�_B�	�ES�&ֶ������p2�m}x4Ŕ�%Ӹ�ib@��8�3��a��I��s��~7a��s�,lN  z� �Mw�-��Kx�+�����PAnG�;m4w��p(׺�zׯ_���7����6q�����Hb����_ę��)T�����#r�;\����}�4���(�>�YN��>� o�՘&�!�>�믪Z���Z�:�Ԏ5f�Y�y�Z�'o=./����x��"^�ʽb���h����7�t���/��=��.㕯z���|�~4̶�K_�&��O���{��~~~7��~7ʕ�-�q��^8s	ϞY\e����}����m6ƀM�!�i���,`椔>�����0H��)�]h%Zu�?|���}A���≸��!2�& ��k^��O-tb�T�sԣR�f��`!�\�N5c�`�dx)O�o�׾��m��0�,;-f��!6���6��nF�^c*� �G�;a5O�=�İ��Z�u����Ђ�RQՑ&�z�^��_A�����2(��"�p�3�>��1Ɉ�Wq.�-r���6�Y�S�[=[�Ej��2�C�`0Hy�
f���PQob�4��d��p����B�l�~��p�m9�g�~����	w�s+~����|���7��_����.a������?�:�	u�\Zp]�EL���w���ġ�,ll����!S��]̼Y��;cH���dLk�N�����;���{�8�n���4��HP�m���\��5AY*r��.	F���>n,���#���~Y�	�fa��r������:h��ʾx`���]PALڇ�}���0
�w<+l���c�[r�_�W?��P���@ܥfIa��ƶ�H�v���n���Ғ������<�i�A>i��/?�u,/�`rnE���S^��'_�7N��kK-�E��)J:��p2��<�^��u�z�X�}�֡�0'�'��[����!���;R���<��a����X���q�f�#�{ei�VG���}ⶣ8rL��/^ē_'O>���	��wQ��w��p�K��3���lӯ,��ҵm��g�EZ��.K૘7lar,�m���J�c�u���
�r���x�׆��f}T-T.������¢c�\�u�°u&7�BSl�a���X(�м)
�O!+0%������ϱغ6��J쵱G5���b\m�"���A�{r�U"U�m	7R�:����v�e��@���oV�CO͑�)?K����h+���iL+L��}=�'�N���E3؎��=W�Д����E$5����_�d�1k���%@�"C8���<ku��	��P�{��ga �d�f�{z��X�i�����'?���� ���9y�ه���l�nv������O|�f���p����4���w?��Z���l��K�Rh�P���y�CS�6�n��>���&KV� �����.+l�f�H���d�;�L��xd䄹��� l��F^��`�A'vQ���_�c�%u�1*�։4��*r/:=.��AX�t3�
���m�N�y�;�(���� ��9�2x�[�pGd���mx���F`4^�ޖ���h�o�oz���������������8x�0�7j�t�*n��>�o>������2>�8�齇P*���s�����װ��T�K(�%�gC.m�\����24,Pqٞ�u-i�ь��6V�iB\ɗ��iW�>��W���}U��61�"Qb[[��S/���ZY��mwZ8q�އ�.���� qhU�2��G�׿�o�vԍ�6~��Z~�t}��b���[@����f�%�ϛ�����J�\��g���h�|�w�Àm_��75T`+���m�,�=�k�N�g)�e��7�R�$@��\��3q��#2���L2���`'0��l�%�.�6����FXϊ_v��zi���禵-��=��0ʹ��?���7VP��^W�҄mbL#lqO(ԛ'�Lz���
,#�]6m���|M�E�L��-�1S�¥�ߌFY1�5����磊��mi��7F#,&��ǅ��'�x)Vu�(�}VIS�A��J}�p���HC��ҕ_)�f5�k��h���U�9���߄�Mv����w����}�%|곏˿7km�L]�K�i	�qcS(|���Kྼ\���ɺ�;ݖ4��)d�8R<�pn�ݤ����� ����.\\�獡�g��V��A�	��/��S����"v�A�j-*�~����|%��p^gŕ����sJu�iB]�|�f�t������c#Ӆ��[>��2ti^Q+�5��h @@����{ģ�w�    IDAT��*_\�s`��4A��A/F��F�B��V��'��.^�*zշ�v�\[̼ZR���O|����Kg1�w�z��P����#wI�v�\���2��+'�Bp��6�9��5<�5�󵅗��٠����	������MbA��E{�G�oa|2��R?�#o׋l�����5�q��*j����/}4Oh��HP.�_�-��s/��۝PH��������137/�G����5|���k�z�*ڡ��;�!��h��)*?"�#
�y�!Ս�A�S�U8�^~�T0�67��ٲ�|_	$,$̔�}sv��:��"��P�F4�G��;�ѿK,�%�m�-=_3�}C�����V'�r8,�����c�ߦ8�2	,e/�^���B�m�)���i�`F�-�b@�?�,��W@�],;~d���zA���.&�6'�:��X��ʴ�[�"d�z(���.ٰ�!Q���C��������c�ȨbP`��2�@?���f,�K,kG��!LCMy��IOyZݭ0��Ѹ���;���G�X���qV,T���16)�9p������~�����	`nwK�	���k��1*{45ioa��ff�x���?-,����h3�]OH5&������),�݅鉲��5�Q ��ғ���A���)Rs�o�rQ�����y���'l��'>�Ad �*wE�2N�
��2ґ�ǰk�5;>�����e3h�
�U���1���
ZH��!�܇�S'�?�z�ზD(���p�q7D������e�Fz�괐/�U�`~��U�� ~����`һf��;N����k�����u��o�<��}�<���������̒���	I�E��-��TT�қK]�x��'ŏ���ƀJ!'V�GM ��DW�Y��/��/����/b{c��[X_���tW�1?��7K����"���59���c��{��	�"}��'_©Spmi) _����X��ƥʴ�ZM� '�[�#fk!�R�6�({D��T�P�|zȢg&3ec�}v0ZS\�Z,-��A��*�/��M�a2^�,���w����#���(�¾0��M�c���,�~�B�ٰX�I[��4�U1b�}R�s[䴉����mm���b#�K8is���@V���j��57�,����H"@�9_J��sw�Hn	1����3�����{zԐw\�VPse�y�-�#��Ye1P����F��vv=���Z3h�6CA\>������Mӏ�p@�,�uen¬W�x6�A�UÏ��;���_���~�-����ϹXټ�CG�JsI�d�􄖄mvi[��~'���$���^�Q�z�]�5����c��`s3��F'N*d��8��?��|׋�/`�L/�_�y�������M�Xf��P^7�@j�;� WΠ�� ��(YԻl���`��-�Lz�f<'���V@��X�����r��AΫ����pr�6R��v�?hca��?}����GQ�Q�ÌQ�R4��9����08N?�:��h�ll�P�T��7��7nl�1^�l�������B���,0W����
^<�����I8�⽲����V�umh�Jm��s�s��H�T�»!�u�Q�eݺ�rdޫ�χ_}T�v?bQs�.��)�����~��,/��'Րt��0M�ݔB";�r�
��������� ��q��O������p��+���q	1|�>�9��=v�2�%bzʕ�Xm.�Ve��!s,�ϊ�à=���'���}�F
�O�h��"�DC}+`dy�|=Ǉ��B,�?[L|x��}��!A��Ɉq���1���f���ߦ��CU��b�C��JNme,�yT0�r�y��'�[������g)� 3Suiaٍ��>�AQ�u@R��|��2^'_��ṬG�d]r��ɓ�h��vWԶ7�^��G�"J!�H������F3f�,Ƴx�̚���q� Fj�7O ��#d�nQmR�)��t�򜤝��p�D:��� ��)Il��xn��ֻ�Ζ�L7�4��R�v=���v�fg����:J��ML�b>+�N;��[�>���?�vD�njZ�����b}��WWpx�$��k���U1�}��"9���9,�l��CZ`^v�Ҹ's���Ɖ�0h�6���`���T%���"	�b[�g���~�2�
'�T�pX�$��m�c��//f*<JL�^�$4�M^�2b��j�P)h�]�� ������b�Uc7̀"M	%�^�]oH���O|Z�ԩ���N/���`�c�:���������'��#�8^��ܼ���uR�x�{R���2���Hz�-��������K��.�&��9g۵�������� ���}w�v-��Mmq�_��u���<�,VWV��h����w61Q,#�aF6@��>T5�i�=~�8�P�k���-(�+�Aa����8������� s�c��ʎ7n����j�U��Vo/���b�b��{cX6P��<h�/Q�����o�!�K�h�sf1#�tPMn�kF�
��K���|�h����V�v�����y4�������K`�s��@:��^�Y�N8���������o����nuJ��:�0�Ӡ��82.�}��,�q��=������g��BY����nm:��J��v��N�#ϕ&���ɻVW�:$͔�B5!��6f<_IF�JŢ��:�m�ҧ7���m�gb9�V.W3D�㗹Ʈ��gM���.xZԷ6KQ+�d��v�RF}B�b�Fy���dU�B��v9Y����q&^T�~��"�/�|�:�r�<9�>�؃��O��ϼ�6<��瑩����/b��G.KSd�����9� -CRmd�kx�p6f	k�T m0�v7�_*����������tj�kS��g��G"���r�����h�0Q�tpx�O�Q����D^�T���pq���
��N��[�i�S�D��I�~�ƀ��A_��O=�I9���:���V76��ɢP��e�!�;7��-����_1�����)����"���������̈́�dˀ�b�EoI��Y[��2�&!:�m��f��.��SB1�qpA������C�V�/��m��3�h��̧����I�������+�{�\*v����)"Q����G�b���8rp�\˫]���\���kXY��G�_A��X�2�0��&���XX��JӐ6H8h��O������e'�pN�Oʪ�_���qٖm�z�*<�u22�
�m����v�1��@�W։LzC3R����Av�۬N,��)��0#R��N�gD��#�2	�Kڞ?jwk��d�e�a�]@�Rg�|�P�7H�dM�c֜9�n�+�+6d�(���SP0����P�@\$x�jxX�a����A��]f�f��.Y9��Ȿ�=�ss�d~0���c�[�@�-�0�cn�f�ܢG� �d��0N��\��as��wS-�����1]�t�2�`�\��ُ�vG\��l����d��#ds
>H�scu7W(��v��c2�(S�CҕĮݮ!먖K�ns7�C!;������`�kVQ�'�Z��I��#�%��w�i���F��@Λd
�&^����w؝�n=�og<t��)z?d)qg����&��&��I��+�F�J�~��$����Ώ&�B�1^"�7��Ĳ%�8| �ï��~�vLV��p�(E�_�xtZ5������������ŋ��_Z^E�u���>
�M��]ss8~�V���G�g�,v/������l����%���K[��:�d)��[ ��ʭ�xp�52��\Do�Ŋ��Є����]�♘�����QLOW17��W��j�g#K���3籾Q�sϟ�7�>���:6�֤���_�bFx�q�[�▃�1�w��݋��ILOM�{X�+�N��+��h��x��.
�[�4��k���~C�V'͔��&(�·
fI���'�Q�#j)�T�=(���{�۲K��+Y�v(�(e�lV	��,Pgj���e���]��N���� p[����"�i&h��Z>ɰ7�9�P.٦�|��&��U�EX &��ٶ١XNu���{��Qsk�69�dp9�x�y�=w�F|���5JdM�g��T/^�ן|��'Dw��q��1TƧ���!��AA������[[2^��fQ*D�L��6�M�����U�lni�i��Y�9�OT5�'Oo��J�1!ކ�'��$��PV�a�N7!��&�����N���4�au/��+U��ɥCUM�o1���q����r�0�u.0�A>��>-agN����5��n6���纾�Kq��s��lP�PM��|M܌>��������%0���c��h+�ҋO-�;v�ıUꤶ�Qji��l�і����w�A��r�8� Ǜ�Z�-?���߅7=���f���<��E"�)@g�zM�lags�N���N~�<����xl�[B��Q�z"EM�7=�t�'N��׼V��"������_bm���`�8��@_1afv�`EA�-�Tj�F?��ظ+�`a�sW <��?�::��Ʈ�2�����q_���Tov�/>!�9{�"�>����ZC�`s�*��8r���(�mr�X���$܇�3��jЭ�����x���k..�d`�"O\�vk�Q/���N8 �;QeՐ�GF�?���n"{*1�"�3�����CU�cJ�[9CyN�5Ľyq�������͠`����g�c�I=bhz����$�C���tT�L>��u|��^�m-V*�h���g
!م_��M��E2D�n�h��{�/���1�B��h�K�==���=�����W���b���ÓO=%4���E�-̋���}{v����д�"�X(wb�k�-^��&Ba��8|�@�d�-�g�� ^>{����rY؎ۇr��b�$,^��j��gk� �Fc�EV��1B\fw!����PI�ך\�$Ri��,���Cvݺ�J�:�E�SL��O�O\(2JP�Q��/ä�&�=���\P[;"kJ.f�:v"�J���5�`�isgmN����-i���`.-�[Z��Yh&3ϰ�xN<h��u����c��!�&���6.�y�p=2I�4@'N�8�Z̉#�s��>���1U)��nt��M��y��߁�fM�Nc���h5�X[_Ş}{����3/��?��O��9{-���j��+���+p��a�~�$}�LW*X� G�A�[�/?���+�aF߯�m�8~� R�@DjH���d���m��i�L{4�^Z��@+���8���~�]����d:腡� ��l��p�ų�=3�O|�sX5���g�?�n���X�شvn9rN�����Sؽ{�4q"���oG�T'����7��ϟ����6[p2:�I�g�G���uF��)�xlgϦ�/|��4��m��IF�t�/3p�?��aY#�%+��A+bc\`2m����i���׭���}h��%����U[�T�i�m/�W�F�^[L�2LlV8\@T��p�E)oL���'�V{-�jK��Ԙ�� ��J�R#�81'��S/��ի����Jw�{��{<�q���4�q�>����_�
D]L�ݏ��TVU.�GG1�tE������c�ZM%�X�zfzZ�R�4�C���Ҳ<��zA�`l��=�g15�� ��t���u�9���F^�BS�yP�OAU4�5
c[g��:@�,�hj�4I���b�(����@���5�s�j�����QOX��c��')��	�E=&oڡ�K���1�QlZ�����}�n�3��,91��o�8l�2c�;@��]G֣!�ڳ��w̎i-W���zd��n�nJ�.�<�[<�)d�F�4�;h�ba9��c����}ѫ�6ph�*+��'���G�'I���Z�m�[ua<���x��\��(����,x�r�	*|��!e<<�WK��;����0Q*c����߇[��������/������CP�����$��g���� m[�9�x�,:r̇�~�)4���tv$�>vXšNߏcGp�p,�om� �{�������]����\���:Z,&%���ɠH�	v/�C������m�k�݃~/�s�)s�����q��
N�#�1���S8��V�������4��}���ő�#3n��2�Z���hǢu��{�@w�i�w,P��*?(^M<O'���J���;��h�{3�[_c�����v�󳟥�P��ָ�V����5����e�(M���	�����$cK��`�&˖�5A[�Z��*�E��hϟ{g/_�Eazl��ݮ��������"ˠ;��+�t����q���
N<V��.��z�zAľ�:���N��j�����bM���:���d��J���6�욝A>�+��kk����[Ȅ�H<����Nc�����h�Tw��(j!���(m]�lv*p+�v�!����}vA�7R�`0�AH��m!3RC[*x�(4Vw��H�e�eƂa���5��/R
f!',BZ1	I�n���3�Z���ݲ@y��r�7%~C8�&��j���O�n�l��	^�A�^�b�.wTd�z�����/�����Y��a��z�7��-G�q��^��'�*�-�,��&V��p���|�"�_����Tp�Z��������^� ��G��c�0QTߞ�=X����LY
.�W��k���_�C��+&?���`F`�`��r��I��D+�����R���Q;�آ��U�2�+�]Sz.��n<���H�^]t3����tO<�v�8w�Eɤ���r�;Q�bQ-�:�7?���}F�'��}ۭx����y#�������'�#�p�6o��3�605�����-��033!0P.�2q�.Zm�|�E$sa�b!3�Q�N�a�i��?�۶�OXFΨ2K �A�ĉ�Q4�O(�7J%0h�w�|n�m�,�L��$f���!8�:����lZ��n�����{��R��e��9~o����k�E�|�h��)N
� �� �>��^<�v���V�=�re\����C�M e��ҵE\�t������\sDC�Hy܄��`�ϕ�U$He[�/zN���r1g�����Ԃ�j[�N411�|���j��NWkD�Y,�#%��A�@wzF�D�l��8�f��D��"�K�n�yV��[�c}��7�D����0� `]�]�*��KDj+���
�P	K�:-��z%_�#v̆(�����B�Đ��Z L\�I91�9@���O��tŒ��F?x��evo�^�
9)���$s/��|�v�>ͷ}ݱ�g�h�1"s?
�3�5�s��'l��S���8�Jt1p05�+���л1��C��#���u�r��n��kx���llb���A[�V]�}�Ad�~����V��[�բJ&��{0i�[�0�/��S��/}�������nEd}G0x��x����1����:x�Si�tQ$C�B-��P,&8�o{�������ov�ꢰ�u��Z���ӧu'�.67�q��%�dj��41L��azzs3s�h���#Gq`�<��+E"V���Ƌ��S�pm���	P��ie�X^N�6��Sӊ����2V���nK�-���{��)H!�9�fP������n6<�*1o�E��@��>���H�[Լ����l)5�|N�8�����TF��/���i���_�X�;嶉���dq�B"�]f+<� �} ll�rT�d�?/�����vq��5�[8��	5������ɋ5,O�Jl��i�L�� �����n:S��p��ޛ��G�*Rcy��1�ژ��=q�/�RX�;T����-�G�WT�04pgQ�^8��!I�B0��Fq/����>-E��Un2q���$�-�c�@3�d���ˤ�TL���\��P`I�]Bʘ8 MP�,ѐ�b`�r1��N��]��3�f��a닡��I͗�/Ĭ�[{��b��
F�h�C�mՐ1I�(Aω��D"��˂�qa�8���#	���G���lV���+C��oߏ�����8�@'q>��ZX[\F�biu/\�,��?�NKhu{�����    IDAT������Ǯ�)=|Xā򾇱r����ϝG��I���Nn��G���y��Y*cB+��P�@#�u�����陌��;璡zN��	p�ݳ�����c{�gv�WGح���µ�:�za�.;� K���U�n�cmm�V( ���� ����6��,�{׻���6#�}�~|䣟�I�ҹ-�1��<z��f4�K��R�1;;�n�"3T*��v���c��Z���p蔮MFC�Z�qf���	��������U�Y���Hc-���$�3Q�v�E:4��6�ϴ�{�i2H[P�`m���u[=l�w	r�3�N�h�0B�A��2p������q�۩iw���ʹ��	9J�͡\���[n�-���.®2 -�+
�5ۘ�܅N��_;^Fx�2��#e��'�p�.J�%U�����Z�y0�����֥bI�Y&"�C����Q�<O&�iڶ�u�������F��P��e��UT�ްsJ��$�>��qؕ݌����=S��
�'�)�d��}Jvn�eb�K�RQ��*/���LބK�Hb���bB$9�V9U��2�$�fjJ2.X�~ό�ϚS7H���p�&�g�4�Q�WQ7χ.;^@	?C�3����Q���f�IJ�f9�s����r��{O�ͯ���.:�6a��%�(�x���Ҫf��v5^� ��Kפ ע�+�b���{�)c����=Ǐ��-�`��'O�ԙeდ����UΚ��"g.K2��0b��(�gW/��+���/e7��G�m��1=�����[v����DlvzR�i�"\Xjb��%��W/�����٨!��P(�;?��)Tշ�(�ʸ���q�q�p����V,���O�*pre\�l�������+%�ģ؎L2?�R)�^��-4�5�e�Y��dWC�ݰ��Iw�vBf�zCЖw��Z'�iRQw}�h��sA��{DqH'���������!�����EE%`��V}O�����|�ѻ� &ʂ&�S7�\���̙T0#�>��(��$Eʄ���B�4x0q�	���o�#�Tؘ�5�6,<�aK|�C@IE���I,�$&�,w���Y$ؘ�Vf����{f��E�F���ͬR's�vTK�@ �CX���$��&.y�F|K:dٹ,�S}an��0�+ۅx����8�����(�1�a̩����q$�b��F�+���$.a�V��XB�.�<)4��y����s{��]��ja��W��
�&��%��:E\��,��&��mI.�z=��	� �,ot6�����	��2�yL��ĮL15����{� !o���+�0����u�'
q,,Lᵯ��dyh�m�kX\����5��,ck�)��v��FW!��W�R���i)��y�'�|T�ed��5�߅\��B��o��_�Ja�wpY��}d��\�%w1p��5��R���,�$dBV�\����r�D��8�u����� �w�����6����0�am��v��l�C�Ur����A�v���ޅRQaf?���'�����s�v}�Wh��4��j�4{�#�.^���
�"ݏ�*eY�d��h&j�0)����۴@4�����,W7�x�}�h��i�ڶ��g4x3�a!�~���-La�+����-'���|����{Cvn�4Y����ʼ��7z�r�
1�u�c$VIPO��j���Q����Œyn���9Q��x��.�=�<}<��3������Gl���J�'K� ���=�礁SY,l�΋������Bθp��AD�υ��c¦A��j�k�=��9j�"Ʀ�B\0��n}&��}G	�m���������(`Ǡ�\�|#��ki�>�l��e)@�SH��\:i��<S��pWE݅ʺ#������nːB�g#Ȟ��r<Z��2�2bi��@��	FH�Z߾_E�0�frݞ.9y_�wb� �711=�~ƃ_���$h��y�{�0If�����i,@�<b�;k�D����{��P��u���16�h��֓�D�Jf���8���u,���j�j�����V099�rUr�8��Ie��8z��-�o<'x�/�c�oF����&���,�YI����Q'زt#'m�0�]����*��&��8�����$h�:{�O����>�vp�B����Z^[�Nc'_P�>��O���LNOh9C�NK�{jbI���ŗ�	���=, .z�S�D�6������L��������� �ζ[���dfN��'_j���S�{�Z�bq�;m}��	���N<�����N[�F����N��ɖ���V(��x�d���Z�zg?��7K�Լ�na��C��m��oad�,�'�'8�q��1~/?�ϴ�;�"�����L��n5����4'��kS�/)0s+O�}����s�-x@�8�<�
�gV�Dk6��E1f���\NE��;M�6M���Ubc2`E�ov�nH�FLqO 'M)l0֚���!/(�$aqD�ײH�hH���@�m_g�+�_>7��Ђ��"�:c�sB��~S5;�*{������]7�Ki�E�n�m
���J�3����@�V]�ϐ�X�~��&m�E���l�����*{e�m�����Q(��w�4�Av�/cb� �L�ϴЍ���\�Q�ڇL&@�ϮͶ|�m>�� m�*�(G"����ƞ�1���G�����~
�MחV�]�%�I�/��f��H+[���ݍb�G�X����&[���e��շ��9-��헞G��J!Axؖ�C��o�U�+d���0�U�GײL��n9�U6ˤ�����Щ�@
]����p��R9>s~��17]G�f'D�ـ����A��Ź/b{g[��'&v��(��Z��P,�ݰ䰴!�K���G}ݵt�:� �U�j.A�9P�(Cg���<��BG��x�HcC��v]6�bݦ͙t&�9�0��k ˴����%{�iC�M��G�#��� n_(\mn�7��v�n���H�p��|�X��s�'��F��LZF�����[�s��ck�$�ԥ���{9�	���yW陎!o��TiM"��Q�2��˩�7F�/=���X�ZY4T+��c5y������(9F��M�0��U� g 	X�fC�����R�Ǩ�W�xV���YڱfkvܸC�g�D%eC�?�.�*��<��"���ә��I2t��p��}��D�M�؆�UeG)�m/[k䏳6����
y[I��p�=$������);�U�~~~��::=E'@?�A�B�:�0l��Q��bl|�(�"`1��F1��%$G������ORwe�(S���	Vf�I��&�n7�������Ⱥ���[��m��-�vjcK����&�_Y¾}���b�����#�C6[Ĺs��ۨV�|n墇͝�8�C��۴�s��(Kk4(�̃Vi<��9v[A()x#Z�f6تL6��"��������pey�t�ce�[��=�
�Kk;��l7BЕcy���&����z���{�`|l7�~Gv�jɔC��E�њ�e�%
`	��SF����WDj����C3�b0u��g}x�MJ��fң��k���ݦ���)yi2�ҕ����p�b��9�Da�Y�̵!���]�u+��;T��3Ӟ�����X�WE{{����A�w��(�bD�_��ÎG�%'#7��e�SM�7yP:�*��84�^�E�s,"�(���Vo�\h->�V�ޜ��â�C	� 1	l� ��K�-�ɝة7G%[P�9�N7��!RŊ�
�mL?x7�a9�g�q�A2�O��_�i�̹v�%������^QPd]A�}�6��i���AtL�>� =Ԁ�ϖ��D*��W|�ct�&z2f�'��� �	�,���7C�kn���"?��e9�61j���K���������Ĳ���RTV��F�6�7:���/"����^G�O �5��J[g����:贸@j�~�н��:�R!��W��
�9���t"d�<���h"i��SSH=#�X@E2y���͍����u������������N�72m�[��%�p���p��YX8���e�LL"컸�H�I���7���a��k�D�e{�]��(�b�d9��d����a�~��0FD�h��m3o	,�P��B`
?�m���M�;,|���&�o�P�;h�Cl5V���k�5�E�A��Z8�Y�;:9z=9'��6�R��v��͢N	L#��Mb4�Ug2�=�K�W-)Vu�3�����M{�4>+�::	T�m���[D�b�5)������D��[e����H'$�9BT�'Ck/��7g���|�N�j[��	^)�rXh��X����5�O�X���x8�D����FL��0�hQ��y>��d�)�oΩe���T�ª�Q��n�IٔB`�E���P�;Ka%�n%4�� �P�j,�b�h��]|�1-�<�����ʄeb:���s� �5��.��#<m��f�n�[�L�B-Z�
EYxL���!!�nD�d�Ф�f�əpM�=��n,)���k�32}�f)�B�#[�/�|��{q�������`'eT[];&�j�[9G��I��۽F}�JL Q���B���ZӨ��p�pb��eL�z�'LMͣ�X�܂��8p+�)U��]hE>&�r*x�I����Fatf��̎)�͠�Ƶ���#�=��u-V�8|`BV�Lv ��s��\E���:3h!��8{qa7A���E���,ң��Pk�`�<�|Η-��^��E*��,cV(�Q*��]�\�T��@qt뫿Ӡ�ŝA;��R/ȳcL?{�\k���Y�I�� D4�9�=��B,��̟Ht�\���
V%]>t��-l����P#�]b�g�@�ac��]���0�����X!��&OH�U#�fg��P�=�Jn�A"Pz�����͸��6ˮ6A��������:�B�%Z�h�ϐ&�@jƦ��x`�)�Y�n;9?ҫlе3Q���&�s�l� ���Q��ٮ�3ь}�(fc�w��u�Q5�o'��<	��O���>�c�d�LDxde'�IqZ�!���2���Y�Ń����$��}��d`b�Q�(�U6Kmg[�}y>��^���dQvI_d���.�"��5ݎ����IUY�� ������ݞw'Q�6{��"�����~�XpA��a�]wZ�P/%�ES݅����;$\�����U��OQG��)#���x]��2�����:v������%�� �����X�c?�>��&����O����<w��\����o<#?��v�:��F�v�Ss'��9$�t�����~_FB�#{ą'ȗ�����O�	:}xh5611�V�&��<| p��S�9;=UE�cj"/����SS4J��=�^��e��汶I��.V�ǵ�+����)�g�FI��QA����Jv���%�Vk�?����)4�Q��M�X���$�&�gԵZ&��z�/_���P4B��C�c��sw��9v/і��E1��!e�.:Y�ݾHi��$G���h1��	mY�]k�:��6;-Kd�g2(��N4w��eÁc�c^x.U�I�k�ͬ������E61>a"����.��CeL�!�j��q3H@��L?��*���vCyڠ`��r��𘂲�<��h�m����+�	 Zi���]���t���3�b�!��T|��d�#�' REA;�UT�.�z�}ن�jX��v-G]�B?�&���>�iѧ���B��ݹ�`����e� �e�����ãQ�����R�LO�>�m��������$F�`�{���{)�b��L�C8��D{��b�f���Y�~���=2=Z�Q����~쳱���_��琶��6�R&����p�	�L�<�U�y�&q�ؗ�@T�"	��t��ڂ,
�>��GE�(K7�kאuK�r�y��kmnb,�o�����|�	
ڠx�-�P�� ����x�cx�[O���r�*�'Peq�	��1��6Q7��|8w��ǉ��(�X5/��Ķm5��q�N	�A�+�%�ʘ`���6�e�NK �����TQh�9n]�F�wH���qu���r͝.:Q�t�`[�1Bf/2x�yj��<"q�aF�� ��'uEm��vV�����xk��g6�|"2�8X������m����PY�"3T����f̹BnRD���b�,��l���E)��������J�"o�6D<�$�F�T��y�����*1���� ���!'�S34����dʫ��w�#�ӄ2���	���g����#�d;i��7R]O��ÌP��Tb�lA��]05p��j�n�`��P��̤LF��a���1e�4�nx�zA��$Y�lɊM��]��G���n�n���Ӭz���6��dD{�Ƴ���o�hL�ź��#b�`v,Z�HY�_n��I�f�����|��/����8�٦>���Ƥ��m���۸ru	g�_��J'�w�m���R3liQ�1�Y�z��\����U� a�f�͟��iqs�8cwL&�F�Hp�H��B]�@4�W��}u�N��5�u%22j`A�C؜ewF�.����/{'�eE���aF�;J@���(����U�;,.-���|��.]�(���&�@��_y��_<����f��|	���'�r�(���Obj�VLN�Fil~��v\E;����Ώ%a��i�],�s"�)Ƨ�~��N����+ak{	S�)2h~N*Ѕ�.za����r���j1u�����o��������L$��8@TfR4①P,�4*�Cx��o-ږhp%�c��Y� ��X�R6%��@:?#^$���Y����������,��^\�X�4�L�x�e���FO�������6�)�'��m��S��_���ai�:��N�j�A������x�mS�Bt�(�E��~���w��QN��r��"�tM`nƼ5a ��g��lf`W����[hS��Xբ��6g�-�F�['%'���m���{u�+�J�7��m�7qY��9��Bҭ������bd=�6�f��Vl�0b#�j�����l�¬��ݎ�<�
�^��&vd�?�R�/����J�291���$�y����
�b40�ش��*��F��ݻ����i0y��y잞���$�Ǫ���Օ�b&�ʸK��3���tv7� �Q�����#��Ҥ�t���Su���S�w6�Ճ1���^��:vn���5;򴪮���������E
��[��r��'EХ����b����A�i�����*�T����鍯���.䲚�m7[���]��4L8�9�(�$��>N�}	��/?';�>}�>�����ݯ|?
���W�}�GDmѧ.��̶��(g��X�-�-�!~;`�!P�g��q��J����h�xRu��R��V��"����
i��j#_��U��+���pĩ���H'��T*����1f�,�&I(����z��fY0x�07������ >�lB̎��᠂����҈�1bR��wayec�*k��o��˹��Xe�:���qH��Xq��Vm��㢧�t�����d�5� &nɒk��|eZ:fo��r���bٮ�D������	ޙs���2�2;9��xdT�5G�V�M�S�̤�]Ƶ���I'4��!�.S�(S�I��c�|簍���:�,��Kc|'<;͌Mӈ}?�]NL{5��n2aa��T�ܒ��|L�r�~1�1���;��-�����{`��{ɸ4��sZT�(��ì���X��N`�G�u�<�]�;]�V���1���=e��)�-r�wH��@B)���?>��!p����Y��B���9�*�"6��15�����xjY�S���vH�C�{�N��7<��R�}�o���pg��^�I\$9�ț۝UZ4���ք�Ġ�����żN����L�Fͩ��+Nzʥ�s0[6hgl�9�*'�42��	mϊ:��zL�5/�A���ĩ�\���[��=��1�x��Θ���_'��q�k�IY=9ip��>�a[*~�"�_^�@�������9�G_��d��@ܝB��B�\�_ΡMe��c2H��)��<��{�a��    IDATnũ��kvNT�8h������0# @�U���})���k1�Y_��\Tj�F����q�zc-b�ҨR����Dv�(��جm�TЛR;����٣�f��a ���P�Xg���o����\B� ��/�)����:�v����%ѷ-�( � &�%��~�c�0��4�E�'ܮ�6rc{�F{��/T���WR�r�ѣCO��0�N`��Q�`��E%v0"d#Qf����mÍ�)C'i�P�ˢ�pj��m��-]n
sp�C#	��BZ�ˍN�h�(g��@����3Z��ĺC�¯��9��"���R���Z�sbpL���σ80'659l�\�a���N»�c=lM������iɜ���BQ��M�+0f̈́�H!w��"�`��x�6���:i�N;�L�V�?sLqX`��gpإiw8���=2?z�ևh��ͅX뤸�����W���%5��$��'�9l����zpI�jkxU��x�� C��W���"I?��̠xE��ETTD�ߟ+H%�0��&Ϝܡ������~����GΜӱ�����k�ce$��IS6�6�Rh���ҟ��`1l�%�&���Ȕ�	��+5��_W��᳜9ᙫ��"466=���l4ٴ�S��U��B����%����=51���#1�p��r��Օ5ƣm��}�O��O)�Y2&������~VI��L�ٽn ��Lx/Q4n����ǫX�l%��s�m�C�����s�mY���C����^*��02�Y����CX,b���H	����6g6.��J�N�n;���˗�k��G��׮���<Q����S�Ľ�{��a�y�}���"����wV�4���킧�}?^x��ҭ�vǬ�R�H��4�%�d.��R�} Cm1��<���tN)�?m�{�Uo�>��g�y�R�~�:���b��92dGOJ�a��7����e��t�.�zTC�N dȇe�u�Z��TB+ކ��!�5$`�`�Z����q8�j�ȅ��`k�����gB�2n��E^u�hu��.����&z*4�y�EIa$u�'�x�.t��K�����l�E�ku���@.�D%�ە�U�I�����2�e��lK���uӀ�n	OQ|�g�����k�2�h_'G�s*�i�A�Ў-�7`� H-env�ͳbR�(����CUu���x1��<��@4Y�f�	3����fx�`����<�۵3{��,4��,J�5��/ޑ�/.e����^���RCOOI2U;�S*��?:���~^j�kB�{�]m͏�?� ��z��v��;���+U5��$"��=�kvk�X��
ݕ�=�wɈ�TI����<��&T�K��6px�j��׬p�a&�c7H�a��P��166$�^{͝�C�+;l��&����f�d�P9Q�
E�HJ6}}*)�*=�%�k��/}�7��ٳwD��\��3��o޴��0,{{3���"<��EhE.z'��`ʔ>{��8�?�ǆ��BW�;H�#�&p�?����.�����}�Z�v����<��ߞ~���O�y�ǰi�~��񾝧�oO���w�	_��Ex���p�EG�>�'��D�6w���#�+��6]!�&�(4΋/��آۙd��.� cY2X��(�?p.^y�5�~��������YS���ob��Y�<y%�1�};n���{�}6nV��5����=��Oƃ�<-M{�^���U�<��?�d}�^�����knG_9���>u����#��M�Q���c��'�_��O(Β!!?O�D%�y�yP�����Ԋ�Y�qP�Q�zV[�e3a(��4�m�AGƤ�����=�݈� F[_Zo@U.��r�;��ݰ	�j6��bqu�:rC�,J���N5i0Ќ���wgp���� ,,"70�����~#y����=TJ���(,Y��Y�d��Q]�?+�����@<l�m��X�ݻɂ��V;�]�Q��8g��O#�P�1�����pty/�����"�A>v.Ѩ�Ј��f���������S��[� �r�u��D����1L�#��X�L�:m��V#��[*�|Edj�+Ɇl]�>ѳI��ڤu�%�6�m��g,��"�#x�Y*]��J��\��c��:� QM�T���j@��.75ޖ��s�9U�#r�,���ٔ�7����xC7��6�e˱r��O3��:�5��#�_+���U���G0k� ~��G�7c&��݄K��q�{�~�h&��W��)�Z�;�8뷏�S眎�O�K�vk�g�w�ސ�r�O�s搖��޹18�y�_�_ܸ�ȗ��20� >��k�v]�)�����Ko[/�X(7�*��a�&B%3�D�r�Gr��^H7�������7��7J_�
s�kضm=��7_t�H}�~ذ8������n�Q�����I-t�������+D����?����_��i|����{��s�x��mC��������=v/��FW�����#+L����8���弼��[X�z܁��J�!��9��hE{n�K�A�X��N�;R9[N�_�X}\}(���G���d�Ҧe$���!��~Ơ�I;%pUʾ�f�J�{�X�ů)nԥ���ц��K�g҆r�ħ� ͺyX�F��%T��[���:똛�]�G�`�hU���Q���������#��a
d�(�!�dF�u������x֍a�.���E!TLk���G����^��D+K2.|�e�1K���͚�]j��M��ܩ�c	*�f�tUL�p*��Fu�:Ւ��0��� Y.��(��I�-��ޘ͠������7���}m��w�������'��$"
�p����'��*R-5"ǫS�R�	z�&&�b�y�p��{���š�m1� �/����dt�bc�PJ�}�f*�{hlrFu©�
��LD,yg^y�m��f����������=��=SN�/�~{���ѡ;�f�o�|噘<]ǈ����'����t�7��|����M �}�d�<�{��}�s���U�;��� ؗ������Ϝ��e���������(V��ENF��q��kЪ5��=c:FG"D�H�w
�~�������j� �
.V�fll�čR
F�������<�w�S��\3�zz�y�q�Y��>��kL&�� �<�s��w�^x;z�,����,�Y�
�?���}ƴ�v���b���� �^V�=�V�n�l��N�SO� ���!�g�M�a�9J�j��'J�+��_
�Ed��jRGF&@�:?a%;I�.%c!'X��5��Pd�Zh��N@�#�4d��aW(V� �a�s�6�W�?��Tggs�c�mή��%sn4����3l}%��l���i Ѕ�H�ķ�� �F������Hor�@?�T��Zf�O7�mlM�Yɸ�?GLv�%�����$��,?��+�ݞ-������9/��dZ�Qt�����s<�30G��ӬD�Mt��A�;�5k����g���}�T\�mt�2�� %��RYC��|�4�5�\�2�&����̗ƴ����YJ$�t����^��&&�|}2�3�8��n�kJ�53�b
fN������ ˉ��6����P7$}m	�����̀��>lx��,�:QCh�d��$A�c��7����8?�����^{G��>{͔�K����8������09tw���}8��#q�a3��|n��6�U���1o�y�����f���ރ{~�2Y֋o|�3����:�cRn��F,I'ǜt.���Y;��na�����??@�����(���z�:m �|�D,_��}�=�baӧNG�2�� ��2��w
K6(b�>�e���$l޼Z~N�����%�`�0O�)�|��j�u��s��'?3h3`�S_����+���(���ux�������������6��_���.�/l���K+p��og�s���d�k� ���X��<���Hztsԋ�Ug�+H#E�p1Q݂��ɈĐ
(�Y�&8�'º'�x#[�4�m�R�R�xH.�r0�l�����}c�]��x�,�>�O����f�ȷ1Y-%.�����������թ8O4�=6了hlЖW��
Lb��%3�(�������i7�H�8��M�Rj�M�B1�{�����v3X���_(��Ȱ�P�T��i���ԗ�%yk�b錦�`ϯJ�wL@�5��A(H(�L�V�X����_����m�A�Y���Дf��="5z���px�� ���q��r�y�!'Z&u��zmفNC�ؔ�C����]c���u�uGi�r��K�����>����ځ �T*��'诔�S�A'����8�:z^,�B���b�H1~��hjIn�I��"�K�K�D���d�D,|s}7=���~3����?#w��G.@�bÚ.8�r�[�3����(
㍺x���ob��o���f�g.>���	xe�J�^t���i=���L��PB��u.ʳ�������+�X��g� w�����j4��
>�����Tq�����Z�;n�8`W��8B��7(�˨���\��>!�����gfK��.&Ɔŉg�;�1o�l�̿��f��vb�8�7��X���+Ls�-���Y�@�F��u�`ɒ�x�u������f����K��O.���������8�1c63�	x^AK�)��>}���/cb(ĜY�����ލ��V~���`��������x=����:��䛘>+�j<N��&�F\���8!��)嘄fÞ�N���R�dY�m~6'RӫOqC��77ِM��My��hNn�+��퓁P�mf�}uwkC"�\����?���e�������h������K�n���I�%���/)5�<�=�mD�)��g�&n,jb���lvĖ�w����m��w��e����w�Z�xw�t��މy<�e&PdcM��r�t[�T���#�3���͎���R�LϏʹ9A�� �<k�����i5�D�]f���v��Ҹ�ѭ��f���6>�����i~:$����D�8;)���b�y�ds����ըWu�'׻TB\�b����R��R��Vr��+v���8}�he��i�b����_�!5O ��R��*R'��c醭����(fS��t��٤��`�>�q�2n���,��g��`7��׷H����?����k�t�����-b��A�u�u2�Xo �q>��Y=�̏ય~T�p.��M0�m+��͔L��s�G~>u�����qn`�.�FZZF�d�_�Y|������W�㸞/���xy�"4j%�8{l��6v��`�U�pr�]ĵ��#��H�q+h�M�i��WbltB\~��8��]A�zf(O�u-����C�ӦO�%�����m'�u�.�Z����!<p��f'�����k�mr��ɓ�������gbx����9䂪��4uo/[�?��,z�U	�}��B-�!'^��!�gNGe�$컯*Ξ5	�=�*��5*�2�p2�:j/Wk��e�E�g��`�d1�SR�+���D=B2oB'
-PP�7��jkf$���X�Z����(}�NV���m��m��e��������g#����Ƀee>O�Äl��ה���|�t��&}=��d�]M�Yc�'34�~���4�d�mL��L>'_�V�]>�Q+�s��|�8ӈ`Z[�Nm�/2��7Qa.�t(�/�G3_jrء�Z��m۷�iǤ�~̜�C7R5$)&�ua�0�5x�X6_��P6/e�6�>N��b�݋'/Б2ɴ����ǳ�6�!�X����3��Ҭ�nG�wA]�Qt��IĊ���)b�9�
(+R��ǦfP���.�Y�#R��L�W�.v�i��8sf3Sn"p�Tw-�!��9�����H�A҈���� -����z��H6��x�5�W93����3���_:U ��kx��G��{o9�3[Y�bۇ6�
'�G���<��\���Zx�o/��.����O��VU�˗��_��N����o� z�E����n��'�7bIg�y#�\��v����ϕ��s��׾�y�g	�X�~n����?��?�����;:QCP,��9H�U���Q��oX��m��g�!FmB��/=w�NpIwX�z_����������wM����=��Wa�:�̃ ��W����8B��'���#��S_����1}�'_�z��xI��_��;�R����y�͜�{�+Vc�@?�t� o2�9���gOԣ݆֭=����yN^���f�*�y�s���ǔI�ؼ��@�fUv
����(�iX65Kcw_�3"Q��M���{�$�Wm<�/ԕ�2�CԀ�L����̖k �Ʀ��d���(Q��b��s�=��Bͮ,��M.���p����Hں"�����9�ƕ�E�xo�.,
�!�u؏��L4](���3�
<���8���DL�J�ғ�b����fa`�q4x�Vj7��n�[,I6� n��D.�\׉j�֬E�X��mC8��E��Z�9�?��Q��n��ڌ�\�V��"��R��{qC���jI�$y�'��VKVwF���h��Y�Hӎ�C>�2v@0�.�vf������*�^��8�����w�E"Wӑ	[��;N=Ǳ�c�˸y v��9�z�������fb����+�:��KRV>hW�^�f�*E��rЗ�(�[K7�!�Ȁ��B�oo��O�oĦ��=��4+�<<�$h�x�G��_�D����8�q�'�.�-��׮�1�Z�a�(B������u�o���˻_���|i�r�g�5N9u.HQ���믾�i�gb�;cx���?����+��@���soĪ����[n�	;�#�y��c�q���F60����8��p��?^ڀj��g`�н$�B4�2�vZ�L�i��hU����E������;��;.����On�	��nÏ|3�0�N��ocɒD�#C��{�
����zmZ��?�]y�eo����}	f�0�g��sl\��`����s�}����W�TRXdή��FY�j;}��Y�_�V�n[�eB/z�E8���fs�l󹇷��+� �(��b@��7;1C�r��#�Bl�J)DeA�&̾y�a"��[������\��6��u����H˚_�m�>~:v�9��yIfkX?�f�l��w��a�q�Qj��ɶ��R0U�H{��"����[��K9��f���C6�nl�fX��Hі���<�$!�~����DU�ؑ�,Ҿ�ynOAx��D�Z7J�#�w���f�r-���
��u�Y�+֭*ؔg��
)��(����:6�]y�0T���L7n�|�"c���ϣ(��E`�&�9��ze��\w�&�K�yM#ϱBT�5����ڕ�FK&�L���W�!�i6�lrU�h�Ii�� �oF4c��fM��������+J9~Os��ci��>:=�v����3sB�6di�\˅So����	<�L��C�olb�6	���J�˵p������N����{~�3y�?��vz����7�r���Q�]r*�8e/��\tϿ�	_��rA�w��f�G�M.�o�������]d|� ��1����I�~����ٴ)Á�g3@���7� �Qu�شx�w�䓯��77��gPvÐ��l�"�2HZ	I$.\�<1q�l�����>u��w��rY�z5�nR���� ��#�n�џ����I�S��5:���~��K���|���q�/E����o�����چ5#���;��.���b�n%T����
s�_�|�l_���x���Ї��#�ƶ1�<�*�&�q��G�BY�"Ƭ)9|�������I8����ҫo�߿�rQ�A��LV�t�͢�M��-����ۺ�%�3�������M�,�u"�F�͘yW㏁�F�<x��u��v����p��Uת�f|�=��L�Neu7������{Z}��A۴A�mV��Kl��9V���1��7    IDAT��l���S`M�=�S��F"�ġ��lV-vx�׀���!e1_*��&)v<��K""PVz��z?��q@�Q�b��Lis�X�l0�&�߭^�[�m���f�r���C��ӦN�V6)YZ���O�1zK��\&	�$mULz!vٖ�2�nK2\ɤ-���"iep�[':��>�u%M���ST)����Q3�i"t�e�C�wW ��Mn���%+�)���%�B9/��G-"t�����4UV�Yh��!��5@3a�q�'`�aǱ��`���0�W[��ax���w���[�yY�ұM��?�r~�#9�����x�O��"X-��M�7�E�iήضX��1|��7���IP�p��C�w
6o*������?�����v�	�􊓔'���������y.s�q`�:���a��u8�S�nn���$̘��mՌ0<q��8N��{�/�u{5�;�(U&�'M��|&�$�Xn$'E�Aս���<�������,����a�`h��V����a��択�w+�?��	��������[s������+��>v�a�8�w�lGm���s�R���i�����E����o�C(�v��Βǽ�ϕ�h������E�V��;b����࠹x��e���Hv[)�8��vѨ��4�h���!�S�e�?�) ����ī���Ə�M��D3�L(�y+E�� R��/�3:k>��5Z�����N�q�?�|t�����z��V�Jm���i�rC��VaH�7��UJ�m�uX1�� �*��-���}"g�`��CWY/gж�=�as�5D�Y8��6��d��ϱ��Jc�V]V�;4@�V.����=:�M���&6�Z����S���P���Sa#��9��T���F�����VQ��8��}}24�����T�;���@K���L��dT�D���q�D|�BOn�(U.s*>�&�n��̂���igz�F�0��
�Gf-Ě�+��4�n4,pL��M]b��Lg(�uR��ҋ���AJs�M�ו�PyשQF��|��@I�^�'��96�J�k�G���%xv�vA���h�����sp���ͅ�cY��\Wu�y����?�zzf W,���. �/ߕ@�}gh+�����~
3wЮ��߀w6P���-�޵�q[����Z�;n��5��/߇�O�kV��&cxH��ٻ���w\�$ތ93�u�yz%��0k��ǧ�³�)�opoD�H�S�M�15�Q?=���5��&&&���Y��?�@��k���?<����c�QM\�'}����Ա��*������|�k���S*8쨝dCz�e�����/��#�/MT�.�~��G>z:x�.��;{-��[x����>����Z[�#pBe�x~�A�50)�A%��(�,�Ej��D�P��ǒM�C���e8H�f�]-�;�6����������c�I3�Z�b��BẔ�j,�8�ϒ�%���3 �[�R ��6�V��hX,�U�S!��4�u*f��4l	�L٘H`6�3}G���&L$��0���0�Xi�����Q�����
�-�n�$#Z2jf�����T<�-�/y��Z�^�IU�M��t��������?Mk�
ȳ)#�Y���s/>��V��c��߳�f:)�������Ҩ�Ok�i!+Q�A�)�:#�l�,���:Ѝ�Of�X��Ce�T���]���#��7ϳ${ڌn�GӍTYMFt��ЌB�|�x>�J��TI�}���a�C�'V���@5Q}�ۃ�?�;����I���0A�r'�#���,[���]��^M�i��,j�X�Ų��X��m��o����"�8�N�%K'6��W����͠�73&��]�8Õ_�/�[�	�׏���`T�P(n��g�3>����V`����7��:*�>���0�"<���*\|ѥ�s�����{��n1w8-׊�A�\\ǅ~��E̜��Ӂiuu��8�C0m�fj۷�x��7��S+���k5k�ꂓ�N�u��ڴᐍ��2�d&yx���
��͋��7�k캳:�S*���a��k�{���5�GPL�Y�Z]���|�����;A�8l��Ф�Ss�}�R�땗��-��y�_�����;��ԏ��>� ��Y�\����{�~T~��������T�z�#8c4��䤸:ʾ~O)�C��&`6V�	Ҥ8���M���#�-G���^N�oV'N��gM-z�ϵ�W1=5&��0�R<�t��̶�Yo�/��t�K�U���x�N��6c�ǵ?�f�º��#�����4�pԊ:�ʘɀx��22Z�4S�0a>P>����M��gk�A����|�//3!*nDHGX;qܩ0�ʧG���
=���93�Ȧ��Jk��몓�z.ا�2��̨R/�if�����=u�4Lh`�I��c��D&�T��@Zg���g}/� d5ђ*�� !0��P{E��q&�@�ڽ=-�{��K%a��'n�t��&k8�	� M��Z����]�Vˤk�F�YJc�ō�X������ݣ4�\�@�M܈	���Z!䀍�D�
�����,�#���7���c��}�E�	�r��R39o��PjRk�z��exs��!���:���(ީxg�Of.$h7j�\���#�^u�ɠ�	3�U����� ��6����;e kV.C��`�YE�y��@���p���|��������sO�>��<���G���߿3g��o�ei��'����/���(�1b`�T$�A����Ͽ�zҔ���w����Cě+'�劢P��A��A��-���B�Y�^|�jGP�׍0>�w��=�=��x��\0�/�3�3����u���H�#[00=��}f��7�%�υs҇�({��;N8ywsn m� ?��1̘6��k8�#dr�k6�Z��]a՜��k1QK�zӧM�P:,�U!ʈ�[��< o4GfMc3��6�'�/#�*�>������bL�j;kt���Ź�,K�r����t�BL4$}����+�ӄ��h_��壕YZ\�~h���	�m*W�)��F�6h���p�?x�)���(�bh�f�@���͍�k�x
��pHƎ����Mb��M6JJ�DA��Rm�-��ՑHX%>�:s�o��"V ���PU�Ʉ����%/Y<T)he���1Z�/�O�Jc<"��C�р+��)J�2*u��16Q��B�Ljs�kJ�~��� E�B2>�6����%"��4�5;��&+:��"�l�6H͒�ec��2I2"d�x�>�����	�k|�����l
�ZO\�1q�n��Ň���(YȦ�Z����|�5�(%��ꫨ!����c����&�mEH�|�h�r��u��4sp3�&�D[����3<��rL��b�V�2\)�U5}B�2d�N�EV݊���8�ԣq�	G���ᜳ�S}ln��A<�������Y}b|%��{/���?o��qG�/~�,]�����y���?N]����;�ܫ0{�=1m���o9K���#lb���p�p���`0�~y<9��FWcpV/n���m7�����;v����G�D�����A��;A%WT��!�\��z����ĉ�҄��7k��k�D���<>Q1d��r,���p�����Q�킴Qr=�4���b��0uvF��]� ��D����-۷��X~�?���-����2~w��8��c�����]C�Th
j6�x�O+q���;�l�@�yhu�a	���pr����W�J���������-%=?~[�P�}�0C¾P�������o�5�S<7�,��b^_����LJ^μ�4��;r�,u��2��۔�Ɍ|U���T4h��`�-L��N�o��zmx1KV����B�뢃X�ܐNx�����k\��&�'W��N]h��U;1:�3K6Ҡ�y����e}�fz"M6h�p�ŞF�H.�`��6���H\W0cW��U�ȋ��//-�����{tY�7wE��M����Y��CC#(Ȩi�V�18��!���޵:�#��_30"B`Y*�2��V��R>�;.NRRB��H��Ve7��3I��خ]���AA��4�X����ϐs�L�9��GIߋ��7k�lD��I++�vnM���qxΰ��Mj�Y��Ж|U�ݦ�'tD�}�*��C��!(�U�do��h������oJ_�ZDm�k��&K����5��d���q��4�-�]�o�܈Ѵ�!WQ�8m`4��N��Oݝ�'"0p��:�}�܋�ʃ?|���}s��S�����D���TxI~��$��v�kKF1������3���[�|P
xA�:�����Ob(�ct�Fv�L����+N�u7>$?���_��ա�ȗv�̝�a��5蟜���M�̹�bۦ<��s���:�v
3v�W�r��`ÀC��h��FK��6��\�Q-]o��Z)&�k���/���?x3f����S�/�=�~s9z���%����3�ϛ�-������ǅg/Ě�U��Q�|_��x���q䁇����^~���0e���y�+x���?�~����>���(Tf���!��U>'A;(;(�9�x�1e�&b�ơ�	a�;*��j��i�:��[�I
"Q� k��T& ɛ6n-��5�vŋM�+_W(����0H�ߨ�`�!�g(����7�L��4'�0u/Rf�֦Nϵ���.����ɘ�.(#�lͶ�}�"�j�<�"ʱ�����C8���M��j.R�+\s�7�Dך��0�~G�T�A��s$2�%h���Ϯ�*��Z�(fH��0��f@�Z�S�At���#9J�{S�"A�K���WAok7nDoY��Ru~h'fe\��vdM�?�e�Fȣ�D��=�<���f���ûf0�>��#��T��PP}|�℗H�k��!�[�T�L-"��iX̬�)�S�c"�n�GD�ė'a�x����aSͬr���l�����~q�)�PSf�!y���d<'A�z3�`;�~��y^[���[���ٳ�a��o/]-C�7ܿ
���c���ז�͍�����ꎏ��Q��l�΂��n������*�>��M��q��s��^xu��Y��Q�?���|I��9���[��G<bc�2�f9�����	?:Pq�0iZ����]������|���N��R_C����c�A���շ�D%�l�J8N"ˑ&��	2�FV8_5�0w���s��KT:��0�mL����2�0}*0w�6=�5�w֏ 0M�����P�"M�F#F���6a˰�3>��{~Ʒ��6�wR661mv͆���ض��*S�Ԇp�e��oϾ��˰��s���wŗ��3DIS����$�9A)D-�0 M�Z�f��)E�X:XЙT���-��<eZE1�j{�%:�9�x�m/���"xu�E�X�����]�� ~Ɣ�;� Á�M&�W}e��#�3^^��K�νM-�c3^�Nm�7��m�dKwt�u.��|
Q
S�k##*�GJ�gDv�O�ҹVXsX���a������a�$Y]l����-���+��8ӡ���&���:��`�2e���r��|1/�һ�D��� ��m�� V�s�	:>QL�e:����>3I��M�|j�:[���H8I�b�I��1�(��7]�a6ͼ�x<��'/�`jt9]�_ CR�5'�P@S���f�f��{2�&3k�k5��u�)��X7W~�Z�6�+�N��|��U)+n�{��닏�&}�R(7�l��L��%S�vP�6�b�F���u�>	ڇ/�/���C�I�����v��k�b{5F═��pS�������z0QA�1���&+��@MO���-h��%5,�{
^_>���i��
�4B�����Qu�D�q������&����0/W@���#��>���bgԡb�>�
���o����DʟRy )bԜ��o��d����x�T�	�.�(���W�U�p�}b^M��������H�����L�Pe*7����#[�y���[ĺ��+��6�p،�PjF/�G��$Y�R)'��SE17�� ����ᥘ<i���Բbf��ۏ���e��,jnC����w�?^^��墿&�8��^���I0c�)�d�V �I�f��ѣ�.FnU�J�j���T�K	Ȼρ�`0�L�Q�����KS�_�LcQ����Z<�V�,�"3i�3hf�4�b~�i���V��>��;�}dpb9.��B��R(�e�n'Ѐ�w�sQ'��(�w������d^�қߗKAd(�Q�T���M(��<t��Z�/� nn�X��<	�U���23�Xf��l�<�1a(_�ϥ�5)h��~�`+Ű�K��qV�
�4sÌ��B���~Y#Amt���$X�>�DR08�/�~|��:ʹ�aU�7ʒR5��\;Gp�67WV	�h'�&�����'��H�S�'�<Ę9}���Ƀ���~#�	~�H��%P搣� ��	���X(�����8C�rx,k��K���S�]�����Y3��4�I74�C�����lW�}�Dr�qA�I%�i4c��B�kj�)D��P#��Ǩ�`��#�WEMFY���eDi��>���Up����7���]op!�~T��\>D3� �����W�Eڌ��3��{X@�P��yR���Uk��U�Y�$��Cr�c���V[(�{�/�q}��L�Vt��#����%ZJ�(�|�$����s9���}��h�}F��9��4���NJd�Pvv~��!�oA�c���8�4j[�3F�6u�U�1��֌�Q��F21����Ȇ���V��X�`dd�|��8&O�!Y���2ĩ�(�@o�T�z����<}yԍ�Z�6�z9�ZJFtJX"pP�&��s���V0�؝k`5��oE��8�0��\7����/G�������=S��E�Crl������VnrB
���ʢ@Z��Qwu��a�Oͤ����D�i���lr��Ǖ&�5b�jl�2`� �i?*�f*�c6�&ǌ&#�}�Z��>N���BSh�2Ej6�e�&l@I��D��_��``F����Q��a�v�k�LOV�؀�_�,�C�%I�=1	�` 7Jn��6�V�`��kMD(���58�R�J�~����f��EW��sSm�
ED��6��ߢ��e�8�IMir���N7���f�e��i	�hZ$b�%�j,�� �U��z��[�#���k�U�v�j娤j�6P���D��� `  �4m��S�kB�L6`n��LTQ��"�*nA�a���T��L���j��Dн��=&��B���l"���k�38h����1�0.#�B�Ƞ>7b�O�4x��i���Qμs')�\N\"f#!�����g�@����������Ρ���N��I�JǕL�!2Nƥ�Y�ˉ�3c��pIk��na��PDE]J�ؕ�C��1�^s�0�[�c0��-���q;�,k��ޛڋg��Z,Q=lݶ�f %�����ĩ�J��KDCBz̊C���GD�8��J|$9�r�RvlT! �G<O�LHS4����hV�"WT��P��Ko�&7���tT(#���Ȋ0��b%�
��VOo~K3�(N��y��%��"8s�!������%_�%v�I9\���\��)�y�]1ˬ��u�r>廘��'�� �6(�I|YF�-GV;�\od���X �h����n��/���\�1�ؚ��"ǖ�`j���x�0#d$=/�1�"�IG"6tLX���j������HLQ4�8��01�Q�X���t�oed�xU��EDxF(��z:y�4@&2����h�heS7�T(����f[t�������y��rJp9D���ᚱ~]�.R��Ko�Ԫ(�Ҭ�ʏMQ��f�f�t��r�1���$�C.c���iI�$S�u��4z3G����sД�b�Lhx�-Bd��X�q��񤊍[��F<Q�[ኦ��4L*������8�v� ��)��h���&N㍚$�\��.ܴt�w��  �IDAT)�2a��K�f��b�-��$��2��fc�)��Cـ�}��%����SOfM!���4���g=I�YC�/?��/f:���8K��)J��J����u*��u��n!%������0W@����!���!|B��
�7C.�Hʡ��z!�_�!�J��W��"qj�`��]�cbp,{�e�$L��g��Oi`��}�X��L�8���Iiī�2U��)`q�@���'�¬*�7Q�h�s�  �A/ϭP�l�_����1��B \���D����f���fF�Wz\fB�af**�/�Km'E$�U�`�JqS��Ά�Qq�7L�5#j�z#�����F�V��ȃ�iGf'|��|lOJ��͝M �"��!�]�Цk�a'*�͆��Lr	��Xs�����TKYr�C��)���~B�p��;	�/�	��YJ�U��D�n|���1���`=����W���r�CfD��0:� U��c=��z��P��D�׬Y� ဓ|O�.Hbe�r]a'>�7j����a�M91�5_�Dm+t��(�͂Um�LEё�0�}�0���ç�;� T%��y̑]���`K�������|?ʦ�X?�jntT�%+f��Yy��M�̯��P�$D���&�f�	MoIy�u��ۍ�b����ՠ:�0�6��/(�wT�:|�7*�1����s��6��s!)A�?�ᱟ ��|i�w�9�ຨgF��CY9_5�2e+1�E]��$�L�b6E�gK]��ԕ�]GS�su�T@VY�LO�f���e�{��P>6�_����3'���UHi���Y|~�:�V����E0MJ)�|�	�;�^�'[2�e:��ԙl��!O�HU2{��@���N&�N�`���ȰMwPn|&��<��6ᑆ�20GRS��/_���!�6/���%�$�����Vf�Y�AHu;���u3�EZ*MeL�#; ��q{Y���li�PM�,n!����v4L�_�*]n��%����Z�@o��!a>�: ��3���"��h������Q�{�&R�Xln<�ժ�G�x���oA�P���R?�1Tkz����Y�,������!#���� �9�A&b�&�� ��$��^�^�ٸE��~"w`�m��#kh\��l��޶Z�؃��J�#��5(�M죈�n�.!�R*(�+��d:s�Cd<�����300J�"��d�,��9���d���W�������GK�~-�(0o�����H���vm+��8F�M���c	S&���'ެ�rY��$�RE9�O�=Q]^�m�%c��b9���ӔX/V�n;tNn�ViOh��zq�gb�8���C��+�x�{���i����:!%W�:��e���K�Y4�}ZI�d�"6j�SC�nb��RSJP�zf�s�_,�9`#w�j�Jڣ�$��Et�/Pk�՞��s�/�䄕4+v1r0Z�BP��r�b�	�����SڙLIk�+7^��N��
c�nl�N.�PK�h���ӏe�:Pa�3�KsIљep��AuTe�L�Z�����`��I!�3+L!�@��C��u�&Z�~1�dT���*%�%�5�5ZhQĥ\F��5SL(���N4*|-������L]�zK{��7%��"d,�eIqj��s�񤮫��+IW�^^7#�!��������k5R�y�C�o����P�Qt��eS�K��|A!�ɗl��O������Zs����% b�����d���L͹``��-�Y6fĝ�E۩��.��NM�U
l)�����Tpt|żҸ���DBI������GH��f�&ם�K�̆�<if��VZ�l7�	M�����"�Ǒgc�X3��/����A�#�䰱9F\�l���L"e0��K�3��H���2kT�T�}Y"%|*��lܼ���-Vc�B��I�|�@=��ET�P]Ha3��|=��$�����Ctl�i��RD ?�S�R�j�2<�6{u�S����=(�ŠxlJss	�)7.f���+rzW��a�9�4��:���1\F�S���e����G�L�G)�FI��H��q��0��L��]����9���'����I�!H\S�(�	'<�S���8L����=�A��$~_�)ۯ�,��*,�Z7�����K�A�V��r�1x��e�U�<WM��7ijÑ�{�Q���r��rF�4[����!�m��ѵ�C��Q�5P*�cR�E)��v٣���}�uN��0uR����Q��
>K�\rR#���e���ȡ����Y�6y�U4ɏ%R�p�?�p�@8	YR��}�!B�}�9
�s)��Q�9f�~;h7�6!�OnsP0*=��&�"���W,HsIpEa��B~��%IAӁ�
r!���0/x)�����&Z4M���8 	P	c�ɕ6b���S9�%43�}�T�c����<Ü�V�on>�g�e�%7�`̰x���Eųiđz݁y#�F�tf$Ҕ%lA&�o����:F2p�)w{�7ޣ�)%�:���rD�ȳr2+�熧���OlJaf�*$D�$�9�0�xB3(B%^'�&Kd��9��6��'!)N�7V3�,�&��q�ĊK�\}n|�yi%ģ�0�M���)A�F:�%��Q,ue0:�NM_�(B|H�P.V��� ��X��פ&/�ZUaY�fVu\��\�
�����s69EGa&fl���D�זO|L�5�a�L�snV�	�F�9�ӄdE�5�d�r��!�K�ޡ*_�Ԅ�J�-Ԩ5�;��:y�օ��lf�q}��+��̀Y=���׼)�E@�#�T_
c�̙Ř�	N&m�81W�l�+�d(#㺹(�Cqd���PJk��uP\���yZ:tUge`/�LLǶ �>i��=a!x�G���|�ށi��fQ!���UPJ��+��hb�B x}���n�Fh,I1} ���F0�8�5���7�(�A���0e��`�Fa*M�z
RC�����yφ7�    IEND�B`�PK   ���X	�O�!N  �U  /   images/32c80dc2-b650-467e-aae3-2893aaf2291b.png컅[K�'����C��0�Kpww ���������-�=w���ܛ�w�}�����鮮���u泒�$**����
��p�DX(��JTTIZT�L��lec#�91I-~'���㇤����4�q���q09���LDq5?iǨ�YÚ1~z��+���g��4�TX�B��a�w��}y�h����v%���&��(�?	�LB�y�T .!>�@�~���c�	³X������0��C����g�t��~�x04ثZ�\�������(��ww�L� �{E����2u���&���ud�	
�M)L��Ok�d;�n:o�H>���ې��|@�X	�����2�d���!+��>P)ܭ��Ș:q��d
F��rQf��}�!~�U��r�AǦ�����mWQ�"�
�f�A������Nv��fj����I�T�b����£*ϑu6��x��b����f:�b�!XAI+�^�guމ3��&�*v�K�D��ϖ/D�Y��,���)kd�V�[��p��H�
L��Kvd8�"���+�0ݳVͿ����C.����S�dV�>Um�E������>��������oHǢ����Jr�ɐ=̎��h��ê��~@'��a�d\Oe���֚�-UWk���c���G#����a&y�δ~S�R�C��O!0����f8�V��ũ�0�S �Z��QD���!LnX��&��0"�^j�4��~�a��p�P�	�����(�T���Sza8P�']�]0�16z��1ND �N�X(M�W����Wb�Ȱ��PCs�_Ӑ������#�z׭��;%,$j�#;�ZH؄�!�eTw�-"H�j: �g7����@��q�'7�����,��V>x���M�G���*Ch��R��N�I%Q&�*WF)��K���#�+��CO.�%�<���K��9�����.�MK�ڂ��IĢsڍ�^�F��<��3��R��>�����#�E\t�$V�jy�rq��}�^
��3i��u$�,c��Y�s �{VS������+��Sr��j�q�o�쬏̝3����Z�F9E�� �0{Q�������ʁ�R.oCq^|&����˄���IFDDDTD�\L�08X���b�̚%F�'�&��ܖ���6�0~9�����'5�ݲD9��[!r������*sϪ=�AsB󣾶$���A�u����ľ��f�+�L2{������x�d!�j�ra�oj�JRʳ�J%��b�,��s�T����ڎ��r�U /��_䅍+����qr��	(�F����фЛ�&�gh(I��T'�'��g��?����w&!^�2@���פU�R�Q�.�Q�P�WY*��z��Q���Z�s���<_2��ֈ�����[�X�KK����V�����j����Jŵ�zysy�!���T<v�Z&��%�Z��Ktֲ�����2Ʊ�����I�I���	�Q�R�ɼ����i�	≉����	�l�т=����,��h�f�dRh��	e)e�1�t�a+fo����'��'��¥ͦRB�YC�����qyp���&-$XM!�S)��i�)[)\)����^'�����ڳ:��j��5j5��j�Jks��Z��&����%�����P{����$�=�湺�˒�֌��e�I���v_����y���|���[��c�,]'_ײ�
�
�
�����j��Nӎ�ܚ�X�z&z~.�SnM���k�Ď�� 0%k�A�nC��H�"�8�:����`�z���9�͙ǯ�5�#�-�M�ڞ�)µ��։����*�YS�KAk���q>�>�>Y7)�?�����>�?D'�2�b�E���Ї��ǀ���G���Y"� Z�0�!r·R�"�k�]�&�sc�2���Q����C��}.�	����|_��{��MK=����s��KB��#�#ԮW���j�)-�wt����& ��,�,�ܰ�2�|n������}���6#O3�����)N�O�I��{!�c�	b�L;�!���4��d|~E��1-�EH�w��D����I�آBa��MH���>�`f^���p��.�R�f�	�j����㩂��U�3����Vemyl��<km�g��s7=���3�:�4�j��:�UA���6ǋ��t�����4�l�>lv2�"������h���oZ'��}���r�i�K�k�>�e3e5�ssz��HR�{����u�nX��؇�K;M�MZ9��ɏ�=K5K!�+Gڵ[^���sZ�Ƶ����ݞ_�^�1�,����<0�Rcc.�l�}{������y7k��>�e����ڛ�츺��8*k[h�H�O�e}Oyu,p��.=�%G�n���O^��ʍ^;Rb�r��
K%;^X)���<�[��m�
c�SY�B���r���%��Q�Q��E��-�p��C�?��­޵g��36�!�	��آ>y��r��S�n��,i��N�-��l[[�����e2pns;lZ�����J��_�ٯ9�?+9��h�o"��[y�v�М�-}�W�δd����{�<\���ж���{������v袀~��{-�Y(Tt7��>�9�,��s��\����C��m��ź�Hm�L�Vd:�Q��\�jrnr|��o�G�/3�.���N6�#M.����ڟ���;��L��B�.��������z}���9�0������Ғ���̏��`	ؗ�zD0��p�QpN�0���R�$��a�^�/�� u�h��-��W	�$9�Ն4����;�AKO{aF��,�~{�Ͱw�����#��$ka�����ňy� f�%������0�0�@8a	�kK�����ӆ���h���̿1��{���AZ8����78�o���w�����Y���������_A�p�AJ���逕V�<��R�rђ��5��e26�71g�u�g~~^�ik�bL�akc���!���@��2����X�ђW"�w2'�d1�������;��yU�$�<|xc�������������d�d������befeez0:{ڹ{0�9S�;��q�̝M��\���Ȟ��ػ��y�Ͽ�Nd�a�?3�9�! ���3�������ʫd�an�-fe��C�������z��������da�ߟ���R���I����"�?�����~�/#��N��f�?|D�g�Of��u��9����Հ3��J�?g�l�,���ä�ީy��/�$��j�=y��j3��	�M�n_L�~���Y2	eaR�;��>,�ȅd�@��ߙ�T�6�2���(�&l����`�yd1��YnP��ܴ����rUV�[/�A}W꽧!�i�[��#����a	�L������Fn�}��*M?���ʶ���__.�SQSK*d�Ӯ�?���0�7Q.ޭU�;R.ELLYw8^�J�����-�4�f9׊O�d����d{���:�]�9h�ջ�T�Qe�\����&	�:���+��FQ+ѐO�~[�SWg� s0_{0�WV)Zhp� נ�Ġ�����aT��M��Q&�t5�܏����+�m�'��i�;��X@!���8ۅ:m^���T#0Ť����\��#�6������JPAv<*g����/��_��7�;�m��w���GsD3�ƃf���)��1��\
�~����A�[�psu��E"2LF8\
4�4�b�ӷ�_����,�J�.!��wg�~�{��X���o�����Kn�O@@7/Fo��>�٧nBM�:�|UtRA=��m�5
հ�d��Ա������1
x�@�3sB�P�?���Q���5݅%DT7Q����b�9�bq`;Y�Lf @�:|bΗ^���| �y�85�֟�-��	��Zh,F2��n��5��o���v|LG��t�WH�.N�(��&�T�ʧ���;��*��jW�ą�ݝ.KsٟU�����*B��uaQ�ޔll���M��\����/�t�݆Ys*���*)!����G˭���*3��y�Y������U_�d��pN�"�^���H2��&�h�6�A��Ւ;��w��QRl,����0��^A^�r��S���p��ܒ��y�l8/jy���Z>�I*��k��j�W��֤�rZ��	E!F
ɨ�m"r��`۟����xgv�����V�g%D9�xTZVd�Q����� ����^S�u�K>����_��^ď}�z��)�p�W���ꌫ�`1���V%��g'/Yn�
M:2�?�#��e�����<\�3�_S�/k4�FU5�ߜ�	~v����qM3�)�V>�G��D����F��㽼��ZFn"��؝*��,���/�jJ��l���!��u�hp��ϰH�\T/�%�V+%e�<+���Gt%�x�v�?7��4����ѠmY��^bx��+Q�`pC���.�4c�8!J$<s����C����]���ܻ��9��.ėP��y���"h3�Ņ��va�g�?����<��#�l4�������ܳ��:�B�,������d���eډvd���J�?��wi(d59�㿟�2��J]1�g����ě/wk�ӆ�q��z5jt���8�E�L0p���(�Y�&���Kia��	�h&�����:��l���f� �2�,����z���}w�k~���G�hۑ�	E���2�2dD�I]�4��g��|oݶ��_5L�"u*��'+��P��o�P��%�0~��Wt��?>�ZO3d�5k�Z'��ϒߜ��'=����5p���`z��_����eƉ+W��h������j�(�ˈ�����U��>[�.��z>��5���mx9ʰ~� ��q�����yE��rpt���˼o�毭��s8�#�좠�8��v<���/	"�K�^��U����3������+	 �V��>s�J������e+���%}+t��;*�-:����Y�Ș-�^���|#�8����и�f��@O/��eo�`���9�D`�hxg�ɦ��K�|���z��z��|MQo�]�~QAf\���=	!����ִ&�N��?S��Ψ5��%+��Jt�ˁ�:h�����ۥ(��r.e6���x���6���[]��u�|��˾�a�#�,A_���������/2l��ͨ W|w�=Ni��[Y[�{��d�$�Rɿ�����it�l��`-/	�����[j��f����E���h3
���)���w�V���笇�y�6��2(/;���#��&]�u�T�*��#a]�)�U'+(�:8>cˈ��ZF6��<��`@��
2�:�3�� Lڎc���������{���u\F|B�QD'm��������,�|��\o$��>^�Ynɇr���{�x�.��CF]��+c��s+9_֎���,�(�$���r����	x��Mt���9�����e/�g�D�v6��C�Gdg��38�5�����`�Sٌ�R���U�Iw"���llT��C��[,\j�|��ތ�l�|�i��jႁ���>\m��g���Z}��?l�����?4t��h��O�'�Z����@~�l	.֪��$�z3dT��5����wh<O6���wl}����:v6}�!�e��摛tKӵ���""A{�##--�Y{ڟ��d�);�%姲9�����T�~�!U�~>�*�16�F^'48��;Z`:�-��M���e0����:���vx	$t�e�v�Wf���+}!k��slq�;qT�Ԃ����"'��\S�T�������"�C�73\���O#Fx�Y����٪���X�B�>tJ<A4n��D:�WnI��
�aV�]�Ȼb0���?5�m��89L��\]$;:}�� �u��TZ'���y��x�ݍd��ޗR��%��Prrv��<O�Z��:��iii��(�ӌ�ް��e�k��fKE�<!J�&ߢ�ى��51w���ĬL�[É���VP�yQ��X�3.~���g���:b{�Ɗ����J�s~�ެ;!��Cџ�H~̵Y�%�<��/�C���(���)��C����_(��iU�Cb;(�>���C�$bמ�9Z���n+�6��"���� ! ���+R-X�,�Ȣ˄���؍#���s�@�i\#qo�W|OO�e����.ċ� �.���.�ق���W�O���[����
>�\v�u�J�c����6KMS䌌�C\�=mf|������uVx[�6�bo���)�U#$CI�!U ���Z�����RV�������^g�r���rXO7$��|t���Ė�l9�NM�|�u����Ə�/������2�N��L��6�R��H<��|P�q`Lԅ��9R�)5
t�4*r�l{�A�.�?K �j9Jf�@��S���I�mi �U��am����w꽞���&&"d�ou�)��?��'�n���_R	s�����y�"E�R2/���(���G�f��
 axY�|�����e_w�����=�
���N ��K%��c�J���>.�šmLؿU��rcd�rU��45�t6*�IT~~;�a�ۢ]������|R%�@�|h��fՀ�B�V>D6⳩M�蒜

�W]���y��\|n�������A�#���IJP�ռ���^�Ɏ0ř�?��ӵ�z����R^	��M9VWyn�^�2�^�V�|���f��Y ��ii���M�0��pZ�?�x��3ƘOn�{��q�.�m�Ct-ۿ��&�*�rl_V�s!���Xp?�@�_����W�>� �_���w���ߋ���q�ɂ��s>��>���0�os q������>�v����aV��w��R�Б|��[-���V@]�Zչ�Ke���l������͙��4��C����r�� x.J9����h5��ɫžl��U,z�i�<�!��D�ǆ�����6��W
���>�%������|��KN��VZZ��[�@�<�g�Q���=��>���N �2�(\�\����ַ�7F����`�f���B��rE�y^Hƀ����k�2��'��]���圣�Rc�̣?<�O��Ƿ0�qX��I����җ����u.E��E�}��$��@�5����P?��E �/�H_}�C.�?����,_�`�gTg��p�5�՜2���\=��D1��#�ȟu�G�OvK*$��� ���;9�7���unY��x^ �9���K�j����Y^�-�C6ѣ��%�%֓[w����;X[��ۑ'[ ܩ�4�l�z�K�t����q���C�C���맷?"a�z��j��L8 �%��Ͳ@ֶV��'�4Ҩ/eLV�B�1�{�iie{�P6Zs�*0��� �?\�'�.%6���Z�o�d��{RL��8�yK����;��^1�_PK�ق{>��'�u����6x��&0�Wt�i�Gl\� %Fzz�eC��5��C�i�5.FXTG
��[����˃��я�V/IbЩ�+��DөsG���q�=%̧�X�j</��?) �:~��2�0KD�ùAz�*�N�,W��!�mN��FS	��uf��-����|��vFs�{�C��S�����M����l�.(����)pߡ`C�P*���R8����U�k����ԃ�Ci�ͼeZ���T��/��M���ߌ�uS2�~��ֺ7�n�si2�i7��˵���%-vCF5���� ~��Hw�O������(
�O�ˇ���q5ɵCu{���>j�2NNJz{�r���>|����w�.:�{�DD���Td�[A�S��Vt�V�3���ɂ�����Gz��u���65���\_,�@��{�[��Z$Io�*l'TA3�����^6��R��K;8x3C��T�.��t�Ak�����<7E�4Ρc��&>����B(`D��QO/���п`;�2�� 1[f$S��w���)X�AJE%�y���'�f�{��~S4M�9�,������c��!�5�@����S�v�Ja�}R���7:hK�qη-��r�Ģ�?�&Z����e����{���s��lSۤ���s��B4-�OB��7w���i�A�kꟋ8� ��Zk��Ǹ��:�]�-ZB��	_
�j��9�B�6dF1�֔��d�=8l˹�<g~�Ny ���Mb��2K;�o-R�eЭ���(�,����,5�˹�������Y�@ޏZ�N�rff�-]#�5q���IX\����H�/V/�i��xz��R�y�B�He�k�9~i�h&;���m����w2<�����*�K���0�<�d~Zt&�Ho<���n���P�p`	�jaW�\�A���B�;�u�$�r2BuCKi�K�DA��Ī�=�#d%�3�P@��26GY�	h�'����� �D�YE��`�����0\r�\�9/w��sA'��b�\qZ�/Z���u�����-��A���p��~����G�y"�:��J4	���� �1C�V��+T�4�'i����e2o6%ܶ��.P��.�&���}0��ϳ!�u�H��c��� �:�t�)��'���M=�(�^Ѕ����?���\�g�S�\|O�t�*Si-���5��ͬ�g�v����]c�Ut
12�ŹȒp|���^��De��э���}p�ھ9Q�Z�K��ދ��$�4��*�n`���V����Z&=A��o�fS&�EU���e����U�Y��A�]d������a���$k鯂tѪrQ�.W0�}�-���<+p�q�Q��`�k��QO�7�����S�*��e�/�Z�5����v�G��%�k�E;�K�#D K���dj��m�$�*��%;��X�>��-]8�*��E-}�q!���~�>�CϗE��hI>VK�l���~�ȃ���:�-t��ySǪڳ}M�,�}�f��:2�W���a�m�����nC8�ȔySnT�s���@{ѫ+C��y�挍���7#z.���=9�{jc�쏯3�8�ؔ	��]ԱpM055=��Q��/p����O���x�(\�k�<��:/��;��i����u�x�S��v��g�{X�Z�c�X|C�9�4��y�}�*���i����mk*o���������f�w���O�K`��M-['T#9����R�x�W�{��>X�kf%�qAgګu��ѐ�W�XHW�b5,,���ݷ�wo)��"N�p���Ф�����.9��־�ϞO��8��s�:a�y��ax#��n�ߋ'9{�����ݐ���>xm�^O�C���-�{���2�0�!5ͻ��LTr��R�m�oPQ�k.鰮e9��a��4n�t�F��&�uk���,��あ|MPJ��a���w?�Ò��R7<Ny�x{y�\���סö׊���]�a����Ҫ
����|()?��Z>l��L���h������{dJ`i�how`�6e�^?�����6I}�%�6N�i5NS�L|8V�����KOV���?��Q{��x�I	���Ԡ�EYc�Q�f�YMt�^�Y���m�d����*G�]R��*�r����ˮ���ęB�n�w��Wm��x�C�&��b{��x�I9�����x�[�yD�)j<t�xy`i��2��3�@�3A�Ȩ��:OBuϗ޵�T��!�3�x�a��F�E|�B�d�NK Փ��q�U 2m!��6q���Żi!>��.��r{��V�o;}o��a�d�q�Lת�n�ІU�َ))�����,����Qe��Uc���,�ݛ����YBR��'�K;}�̏s[��I-�ک�}/}��N�������0�/+�y:�n���cc:˭�X�ZX�d�/��(yNJb>g�6�A�P8���!bb�t�~R|rc(sq�}U�U~;�aP�W��;ǲ��bo���nZ��p�������ͱ=���v��|���Q1��D6M���ʱ44⥐=q�,/k��&�	D^i���rW�ڑ�VV(�K�H���v?!�lx4��}4^k|��6x˟���s�b�6T�� B�DJ��r7���P7?�S��αW-��`���R񞷒�I'��s#���DS���/BʦN��*lj�X[�gn�C]����m,��&4��1��=غ$B�^�ˏ7[��Ǎ�O]���o{��}Ҵ\��ZsE�������g�A��Visd�b=��XJm�"��u?&*^����C��"�zqہw*s˕���N�$�'�{�K�͵���PS���U�[��zˇU�,��5�ĨU4��y�n*��[K�J�.�쐶&�v.U�H�W���x���1&m['6l1������q~�Ho/u��^s
6'Ն������"����[�<��:rw�p�R%��9]�����N�.�g��(��m�/���|W��^��;�ȵ�w+� A�"�o�YN���>#���i$o�2�B�!��|]���ll�.��)D6ەy]�&���:��N��3�c��o�t�g��b���&�/�ڵ�%'������5pq���_�l�C����f����]����6�]�3�ܜg�XԬ����<�K�0�N��.�xxMY��bUW�AI�|���8XxK��c���ǆ#C1U��]ssU,K�UkA�u�焴IZMF�W���|�Q�3w+~V���35��x�|��o4�:���PiP�����x]؃�'<������ٔ���m�y��DU<x����Z�}�Nz���?��c�Mf��� �؞�[ȏ4y';�-�4�`��������?~��5"���$I��=���a��:�`��sd.�ڋG��V¦z��o��Śb�p��>
��^��]�PE�zi�O}gj�8d������@p�m�r��+t�B�װʐ��^�eg����2�ݡ�u�AW���}6N�KNO���{��;P�S���~�'�:�p�0ItbH����j��@��`M��3��*�]Eg�~�qtA�	��4��9s#Z���+W���z�`@L�q�*1_F�����l���3hT٩�����1dp};�(]���"��|l+s�֖�n�ң��P�N%�@�_�V�� LM�yC) K�v���N����3����
��F��3�_�D
 Q�u�e��D`kUյ�zt�{������(g[����~M�=����C���P4�IU��*2x���Oh������`�H��"���UJ(G�~o�W	�D����,{P�pٌS���F<��Z+��;�U=0i�1��2�U^�P#�1`���wZ��wZ�|�A���aMv��i��47�]�j^N��nM����h��v���u�%@��h:�#���z�t���5s����6S�.ח7�� װ&p'� �=�+#��K�Ӓ9R��������H�	9����I̙D��L ���B�����F)�1T�����.����6�	og�¹u��IDΘ�Zn�.^rl�pG�[e�DN/�@��4w#H�\���G����}�˞1rb�`}��F|V��e��Ev%�M!N����?Zd�z�F�ֿv~^����)�z9��^�+��=����$�͵4�>.9#��.����1����B��*�`�3[~���%�:t{��kU'<ǘ�l�8t�]Ͱ]�b�&y5!��8֤U�U���,R��ά.�w��+�ѭW:�X�W�-3B�G{�#g:���N��Ew&�a�ߨ����\������e	3Mۆ�ٻ/(V��<۹^H�Tٽ�I�%�FCߨ���UV!��JwVOh���4�~���F~�S�`{�c�Q����P_�ș}�.��؛q��;����݄���a�ؙ�\����-�E'Äk,n݀�E���lD����i�����*��9PC�/j0rÃ��I��;�JX}�jUٶ���L��͜OAss��ϾP˜�"|�n��6[��4ʰ,�9��I8�[��a-�7s�o��\?��z�#Q�y����3�{Oaй��!���GZ {/[|��i9)�:��Ku�:�l��jg����?
Hk�w��|� ��
8�$�"��[��`��p��`EZ�ޅ����h�X�R>��z�\�`�*����ń���]��R����^<nך[�I��-As���(��m_OIF��n���m;u�و�3Ξ�
��}��ߣA�[���D���{Y�;�<�n�,��[+�~p��x��;ߎi@��_$���j�h�ߍ{�%u�qx(^�e�En����f��6n������_�E�v�{y��_Ul���d�:����$��d��m���` �p���P\���ŮTVX��UyN�|�+� �K��@
��"�O�ɟ���6�ME�Lg��厛)��SU�՘���k���1\��s�~ߪBCi��A|��\qZO�"q�t��X9�|M���K�=н��a�c�^[iO)�TT�|���Ү�<��Cj����c^�i �)��Q���Na!گ��E�r60x�a����������FqM�ݏL=�ʜ� l�6r2e��xd�Q�WP��̽Ӫ@y��?9��y�thg}�3bj&F\?���I6�!_��*���[�,W`�]�+&�uU!!`�s�{jv�ܩ�����D�z�:�#E|fzB:	-%�_����G�#G�c�|G������dd1�Sb���z� ����3.Hh����FWwR*�<T܆!5v��j{Ӻ��k�L6׽s�M#�%��쮪�>�=���A��[�ڌ �|A�"E��-�7{��n��M�DKu�.�!�!�+�S�������?��3Yy��p���<��p�f�{�@�s�蝎�O*-�O[�Cm�?m�-_���j�Z�$�=:��IhO���s���d~�'�d�?#��1�(�ɬaA��}{s�����F'|����(�ʣ]'p[8G������M�	Ln#��b��en�4my�@@·�0�0!�������mE��](���5 ��i�(��v��@F�V?���8ݬ27�';�%x�D�;�ݡ���ŝ�M�3c?+�b�=�ͳM_�o�����P\b����w\؟����VWG2d��[:0���,_ v�����`�a��tP3�;g��t��k�ޙ�m�EQl�����F2�"	/MV]�u�o)�)1��V�ȣ#�k�fy�����0�-��3���4u��R��>����9֫6c�(�Zc/0�O���G��<j���u�Q~��]Ȏ�!I�YJ��nU����+AD���l}7����M�p�����(.Y)S�bs<���>j@�ք�������P��*)IA����4��S��8�$������s��5Գya���@�j_���&���~��:�+D�5T��JU`h���-��� ���R�c���m��}�I��Y��W�݅��" ����&Nq�j_8���Cqk�����q�o;�_�29s�Q�Y�)1�ݖ��{���:��
&y��
k�>hs�6�<v9ϱ�a��v�G���|�5�( ��ZH"�<���@|[�OѰH�&+�m�
u�A�9oD�c_�K3��~'��h�f2�v�ŕ>w��p�>�4�э��]<��b�#~��N�֮��V����1O�Wd��� /`��M�X�Ȉ#�;�+����k���O�h����ֳ�E�ռ�th/]8����A%��c��|�N,�Z#�e634��M��W.j�ȏ�{�
7"��wX2S,	
k(�[�QX�d;N^@�N���=rr�5|����V9�L�S�~ߣ�q�����d7���Õ8����ׇn�k�H��(3�?I������oO��߮;.��k,Ҷn��
uED+٘�翶[|a��8��A��3����~�[���쁽�]�ן��=�a�2����>&8�����\��6CW��֕�R��J.ܯ}�r=�����[уZ����L��G�ڶA����(�a���8����U���>��Y��v���I�}F��Ji�p}��0��NXe/��q ,��ܲ���b�f���(�ǽHv�Tr�92oq�i���C�I���_�0��qE�E����>�5�{�3�������P��{��%���ϫ쌓kb�#�?�4���mMȦ__|kD-y��ީP�M�ƃ�!TC9fd�8d�q�Y����)��cDu�A�ٚ����=�U'�LC�)w�;q;��E�Ť��^��(�v;|�����Q����-�h�^�
��d�8�TN��R;�Eo���P��1^A�(9��V�m+ņĕ�mf<����\ŭ���	x͇VD��(/`%M�䒟�R'�p�C`�%��Ü�2c�bm�*y;�Mi����S��H�p��W*��} �^�\�Trt�Q&3�7��NVHݹ��nHx�N���NJkp��Z��j��߉�xÄ)k�:7i�]��L<�k��6󽭋�>�v%�j6�y��ks��S�y��׵�EJ�@�/���5��e��y�~|L���cY�i��������Ԃ}Y�y����V�#�]Kɕզ��޸��A�ව,���)�A������Rz�*�%2��.+��
����]�*��-�<mkHs���s���Bra?D@�8S��mm�[C�p뫪W�C�+zVX�%6�ԌF���Ү���pȔe���b���0�,�w��w	�MH@���B�T���|c���%9��� ��f�0�8 [��`%B��R�8�А�
�_Hl+'�h@W)���DH�S���!�i�����
�����I���1���jV/`{�a�ܥ����� ���� �� <�
��2YL 73���``Paا�A���c��t�����OO;{� ����@�@�����g@��pq� ���Ld!>}����A �-�˧�Q��<�1���Oe(��SM��Ӧ'n� �0�y�8G�����Q <㉦�"h������� ��iӈ=U������C�XS�i�y��s{����j�PF�E���V��$�-�0��D�'��
Е�~K�o�v g���=S��W+�M
,OU�.*2�	��L����/�a%��ug�?b⎉v}{�ߚ���׌����`�I'.e�7]�����~��T=!iPi"^��%��rTx||<N�k���ĺ�h)5�}����T��#��<d)� [�;0O6y`�����Ww\|��o�S�����vm����Jӎ&Ým�:�>۪�/X�vR����%����l�Dy�O�l�!�ŴGJCC#�i<W_Ч��`�Vi�כ � ���jM�w���Sٔ#^�ñT������;$�OI�vv��$�Z˞[ĺnc_$�<O��88��.M�>}	��,}u�����x��MID?�~��q6u@J,J��j3Wa؞��е���W��������(��G�rK�i�~� ��S�n�D�G
k\�e�W|,�w����n{�C�}ǭjE*����E���je:S�~+m�U惸ڵ���=ǿE�w�]���ϯN�u];�3�����4rXBG�k|�H����Qxh@&m�� =#RZf&�3t��8*���	%N�e�^�b308uz�{��7�p:� �`P����5��e�+�r�kA��������l_eP�0��,�N�X�N&{�68�}��\NC������u)�\x7�֫��X;�q���N��V�_�Ss-�X�W =�_.w��ڑK�͵���]a��B�	��VoO�z_%m&r���$R0�y9��n���i�'�!|r���d&�r�xL��	d+#��z�5�s	.�S�Tʤ:���e�H�z�a��ve'�ow3��Mv;~h��|kU���5e1L�����/+�.��ӿ՞,��f1�C�|?�f�U4�X��}�;�0E|�g4�E�i��KJ>)�%���vM��	�׋�̡S��oG�g�]��us%�̏&�B�1�N9�z����ԳPX�S�-��p��FW�s2�,����[W\KmSA�s�Xl����w~P��[_z����ط��R��t���w.���Ӱ�y�"�e��\z�Vt�=9��V�O�A�`>�|��V����/�/�!���;P�{��x$,nԸ�J	7�R=�T́�٨MKxXI��� ��v�H�Ϸ�>�������(��Tg��EY3�\S�^�:�;աSn�L��pi*��{m�P�4�����#�2��ߊ�S�uhÁM%�X�-���l7.`�gl!�Ov��svW��P?��UWmRq^R9aC:A�>���H�	��o���MG�ߝ��ُ��m�Nd�QڀT�ZKS�G�7k��ϑ`��h�_�݀A��ෟ��p��7Dp�D�Zz��-��P�_�F[*Hⳕ�6�$���L�b���O<���"`#K0����i`i%2�������1cy��OU�.S�4xKl"�5l�[/3��+�.�U[��(�sbX�y�L��S+^�P$��r�^���8��-����H�"#$��]�Nz2�耣�(���]xV��ȶ��}�%�����0��u�}��#g_��\��f�09�lE][�����tm���_�O?���sg:�����^���1��0_�ؐntڀ0�>�Y����<:�֮v�&:y���Tq�F�~����'tZ��w�V��K�6S��CՀf̸E�Lʙ��uM���x>�29�9�$�,a���B�ҌܦK���źQ��Z8Ж���V��t�tFh�">�%�$��c���[�NY0<7�'�1@_��Sr�4�n��ݾ��������D�_�I��X�&mD��|�U��dfC���4/�%�p\F��T�W*���KM������ע+!s�s��������0h�/�J!�x	���r����%S�0#!6��I0�Wף��>�`23�%\f��oi�0�)�y��c�Zϔg@�y�G-��崳}�D��I��W9g�u���[�ŭۍ�h�l�����&e��ɾ�-K����FQ�2-!�fO=J�%31�"�0Ӎ15��;Ռ��z������s]��y����O��$V�{/)6��&ڷ����n�n``����?���e�fI��h����Y�)30"�r���,��[w@�0���S���;ƏZ?��7��ߟ�?�m{�۳��/�R�~f,�A��q���v���M{�5m|�	�j7����No�X_�*�]�2� �Ш�$��*]�����bQ|���o�#mUrVk+�k$E#X��[a P��BwH�����d�~#F�_?�y�{���.���G��9s�4�/��x6a5K\�أ5f����ǎ�ݚ����_ ��T;|�,s]V[�jO���Y¥�J}��H��U� b�u�ڽ�:&�ii��^B�x��ܓ&]z"]~�`����&
�Y�[�Y�I."ql���� \ô����Z+�ˑ:0����J�}�g�y�A�v*��E3�����!s�������.}W����&��d3�D�}K
�y�)�
x�m�&�!}1��t�����E�křҙ�Ww�Nާ���u�᱁�O�L!$������B��A�C$ ���mP���i��Tm��s�ǐ�6޴{ �X�$n}Oni�B�9�]��:��7��+�ݛ�p�]����^F����j5ӂ&�R;;�F���	��/�sl�x��#O���,�&��
i�?���!c2�(��Þ���.o�@��DC�HWb���Lż�ӱAo��m�0�~+UJU�O�9�Ȓc�k$�J5��HF��pT��؀�Ǘ��$ ��/�w����/�yʎ�a���6iI��⺌��C��MY��n����^�����1Jhc^��r@���I�L^7��!Ebddd	��(�����,�������f�"/�����s3�$�5�j�������� ���@����A�O/��iv~���Mr#�L�2�������"���|�m�K�����v�yTv��>`h��S��V�L�U~{�FB?rF��Aq���lT����������uyh`�mG�OS�*P���9d]�	���@����9��-�ڂ��[X��.E�rn��<��L-6��͠��7}@:��op��W�z!�Kv� Tꓴܛ,�����	�J�r�Z�	L���u���ʌ��h9��s�*xp�6P,�uqo�o�`J{˽G�:��t�lq���Rg��#~3d����m:��:�ٱ�b��(�����ع��WB�(@��>?�Y����-�����D��Ð���`����D�����H����cmO�4���� T�3�[`�8DE�b�>�����Hu�0�f�^�럶 �����z��ϻr���qKrXs�S~x
�i���V��]��My��E�C��2&/�ܣ�mn
כ�\q����ɽu�A:����u�p	��&
Ό3Ep:�Y�-Z��z#�4S�
#�0w�z@���R1�ʥ����/�j1@��wlf���{��� �3����""�by�2R���Lu�?��G��"Ȭ[J&Ɓ��nd�p����3��?7SXq�%�b�'��+<2� �/��z�,�-ڱn�ԅ)��>e�́��sOP�Xiy���{�Fi��58�32*
A�*̒�&�:$'�X��M��H�Y5���73x�!�]\���UŖ(�Z�I9�Lw�C��j'�>�(��c[t~e�
��I�3΢&E ��k����qRV�7Z.������jrZ/�R�OYv#�I"�;{������۫$��KaH�k+��aS������Jl�R��ElxA�^�B��/{�?c>s�#���`ѧ�����#��/�;�5r����k�Ik8�4�:�gC���MH�JJ����y�%�Bya�oB�"�^P}�H�x�b�?��<�b�aOå�q^ƹ����@�\��U�{7�F^�˃��Ҟ�w��8�x!d��v�ň��f��%Ɔ�h���P��l��ss����ľl-��K+��p�d�~+
�
H|\���	�����8oC�y�k�e�.Q�)�z��D�(��M��Ғ�'�24r�G\f��"������o�pq��P���>��܂�Wt��招��'3$΋����-�6�y�x�Vǻ��Ҁ��?��s�J+T����f�~���A��O�J�]���Yi�	�kdw��x][�}�D&%��c������I (�'W��31'�\Z���i���Wǀ�B-Po�5�V؜#�^���
jUr��� �3A�KI,_k.�h���&E��������˦;P rn��|qƤ���z?��k9u
����Dʡ��%6k���w��M�»����`&�6]i2^��H�qm��W��l7�]�yq�f�3��}�f��ϟ�eھ�5��	�hy\�/}ePs�|�0����_���T��u���櫚!^��.O�^$WD��bm�ov�֓y��
�y� 2Wr=$��B�C>Ƨ?[Kl[Y���� �s"\@�����!�I�rȝ��n_UB�������.�]sa��V��E59h�����)+60ߓ��<k�+�FZOn��w�2�Ckι�[�>�O�����y��i��R�w3�{�җ�Ϋ����d|@��0�Ǖ��7�y
;�i��ҙ�-
��y�x$�jQ���z�� �l&޳�2�͡A���b(�l��������`DM�@�Y�a�⥩���q���c��H�ڌ�>�M��1}V��`!�C1�ݽ�3S�\+¼�|��8:a	6'�Ƴ�n��v���3;��KM�Co��W�_��	��6�z���D�O��پ����J)�{��6O��vRN85b!�y l����e�[g�~���7�oyl�y������G�>I�PK   ���Xp�֣m	  (  /   images/37476977-ab57-4ec9-9e81-825006455165.png�V}\����:!����/	���l��#ɤTJk�×�)���KS��L[[�����>7?�V73M���w����ͷM�f�/���>�m�������{�s�����<�|l�؂Z�� +�	A�I �!���'��	��[A���cEz��c�h��}��{0$8�0���˒_f� G@���#��~;[@p�b�I�X�����kk�̒%$#*��sTB*�+�Kj{A�������0Z�0���0�K�$%/`$4 &q�q8IR�@D�<h@6�)܂���@Bt�v\�0���@����2���Z$3d	V���bq2�BIOO'�H��(�����:ʺu^��K�!�I��ՋA��arE	��d1_(���q��C�@a�g�Y܈+����@�t,p@��B�&S)��6�7ki��n�n&?	��A��_@�K�_"���P�DF�o�.75X��b��7����m"(��b�)Ky�/��vg�e���A"��d�T���
\:�=Y[b��y�=7��.�_U�f��QՅ������cp�-��8X��|.>;��7�����k(�'����5��2mZ0�>�V7� ž�t��0b(t���1�s-��[���J�K~U�����	z��
):_���F'4Y��>�W)6o����=/�-�dX�D����G����N��l}g��1��A��$�g�D�T������-~3�::�̰�rϲ)bP�ҽ6]RҦmh/�_j�%�'fgn|�m�YAҷ��I*[�^d�7�����\�g�;[�=�������~�U�-VֳJ�C���Y৺ҹ~ �^�Z��p�w%�F�z���=��h�H�p�O�{��O��j�K	�2ӗ�U)�K8-f�;(y�'a��s��V�-*|+�#n�}��:+AF\R�w�~��0+.ɕg��r�-y���|o�Z�,�߇�$�V�,�0�K�p��^�?	p�T3NB��L?����mل6z�v�����~�S��|>�S����1�����YX���ݻ��Ϗ��޾+:����M"7ZP�n�;����%��ae��I�s�sָ���p��
�(u�h�M�Vr\>�E[���p�֮GA{�E�n�;J�e�z�6Du{�����LnR��w�,�"
��|-<*s�V��Ի���}�ބR%��u=�șk
r,9ֽRf
��E hc�$Q�U�b?������*yw���c��k(U����N���y���#
�G '� wF�/H	2c����=���O���oƊW�]�6���٦�(�'D�3؅���|6Ex��J��t��4v�}���ʰep���z�E��J[p��?6^o��k��<�CH+���]j�@,^]�lp��i�筪�
R�q�Bj���!�A���TG{㝸lx�z)]��%�T�-?-;�9̂eF&����O"g����F('�p��`��-Wd&ܚR$l-�4�ND���]]�+��{�]]�y&�O�as��%��z<�6j��	��CŹ
��p)B"h���K���:|)e���'�ܮhmU���׮�g����颏�B`%�(���3��@���&�4�=0�5�5�z�x8e���mE�k�_^�?CR>���$V8��s"q}ֳ��c�y�-����go ���� �z"�1���t�����"����%3�M
����6~�	�����X:�Gc��>���sr7cS�I��ʜz虙9>�#���vt��h��q���=ņ��3�(��)�u�l���p���DI�.��=��XY� =���]k��lN��i�;��_�f�[E0�������A�S͞�Wl��f�^#qbȰ��}o/Gh��Q�l'֗�"�M �P!|«��ug�{�@��9��:�oU?A��0�v~s��Ѻfx��^Wz�27�лW��9)�ܼ�����X9%�+�O����R�c�v5n`XǦ�HI�=
Xĥ��I���t�~�ș4�Tfv��V��jtCV�g��3���<~x�J0!��@�v�髙 ��ǜϞ>{8����4�}��?�r������2��E�+@ӢS�Kl2�]C�U� :�gg�S3�v�.U��a�WV����#�I8gϞ݃�)�$Km�a�gr���㏤��f�!韃��9ho�B�uH���y.*^������~[Տpfw�fu����x��P�dTq�n���6��>%PF����YQk79H�.e�C�B��<���է���-��G�qM����(I��ވLx����Bw�crQ����uK6�U�_)9�~���F�d���ΐ�zv|tϧ/��g�-&�X���AE��K��JՍN�T�ᬇSo&4��}N��;���=��0��W>A$oP�����B�,OxbjM�`�������+�PK   ���Xf1:Ϫ�  ��  /   images/385d3502-8778-4b9c-b5b1-c060638a35dd.png��eT\A�.���;ww��{pwgp���tp� ���!���;�}�sκ��w/��ڻ�������Z�-EL424Le%9�*�]���"��-}�z*���1�ް�:�Џ�vF���ʬ0(�fXxX(��`�ђЛ����v�G�Gk���b$����?Ox���H����������e"��A��r���*+C��6�vv�>���1y��'=#_#u5Q7N+[k;� 7�<��P���׊&����G4@���Q(�������_	:#u-Yo;ANnNn:I4qo[{Q9���C�$�}}=E��   '����ہ�GDD�������:��'���*��݇�?B�G�����������;�뻕����������"� ������fA�z������_�_ſ~�r
�s5�sr���C��WP���:��4�?9��ON��oN};oY7谯���������q����q3��,�&���b&�&r��3z�,'�P|և�kg(�9jr]�4z܇��� ([��̩��u��#D������p�/�2�(((� zy�^�$��%`�I{�#��#~�28�*g^��>�F;�����(�6Fͳj0�(
\.'�&Q����n��u��8c6a�k�����'x��a��q�B=�V��k߷3�O�KT`�e��RX��ꀌ�����9J{5ډ�?�l2������_�	^`�N�~�����dɍ���f�h!Uv,�3��øӓN�6 ]Ͷ����}����b��q��&�;o�x\A�"�.��~���#�W���Un�l���(޴/��\x"�\��yf�Z�&�ά������Pْ��/�����d��gRїAͦ��>W�7?�j�����\�
΄
.�B�K]ө�Zp�Q�T���\��w#)L5����ILqKDX8����$YN�?@9�o���:>A�(��%/]�j�a���$:Z6pnk�P�A�f[�~�*T�����5x�O{�4���ڏDWCR�J�iޜ$i���E3�f<��Ӌ��!~]%�܂�4\�����;;��L�����bvԽ��J^�����`�4���˳��s���VM���^�O���ڦ��ee�����.��O=K�~������h�J�e黝�զ�����C�� ��������F�����I8M��%�y��^�$|�xht����m���]�e@(�8�;��ޤv�Lx�}���i�I�*���ò)�>����-��د[�T���|<=\?G@���f&��7��տ{�/����0)��@��1����xt�Y�J�8��FY-~���
�s�?,\�y���:?a�d�C��SMpޏ�{Mw@L�#N/�i��iâB6��o/1�V�C�0;�Wwx���]�l�l�h<����A"����P��0���?~�˖�Tm�j��B4���ƨ
�^�tS����\&�a(���:��`�����~ȁ�@0'�����@��-M�v��j�s�u�D&��0t���Vl���T.��Â�~�6�^]��Z�C�.ܬ�+������?����|7~�%�7*AX�
鏖��u�P�aY�:DkvÝ�09l���Is��p�oH5|��.��S������a��I>G�S�j��p=}T���d�t* &����3I||�Y�U:L*��)�B<%~\�ٹT�B�^� �^&k�/̟����+M����&�
�h����*
�>�)�׋�]��7���Z
(�y���(7�=�*��tQ�I*Q
3(��[8jx�l��.��lJ�(\8�hܴo!�;|UˀKP���;�&�#�����4{hf��8��b��@�a稌A��	��'S������\R1�k��C͆-���\N�f�Z�f�?Bv��g�Ͻ�� ��ӻ'r�5^����?��6��h"W�\E�d9Т�良�W��@o.�3��������I�>k��8q`�A�{k��<V���k�߿ �nC���c|�9�l<�;'��D��8�F��3GA>��N���^�
���R�n��ہf!V��������W�4�'��3���v�2�-愤����Z�V�>���?9���q)���Ӳ p,5����ɝP�q¹���/5�N��l� ������J����� �Ⱌ :�Z�c!��f��rӼ��0{�a/��Ӧ�D�
�8�f�<�;�����"N�Ě@Ϗ�FD;*��y}t�x�������7�/��LY�z�)Hi
}3�z<��Vϯ��azrg��q�aa�.�B�3�$w��#Û�ÅSߪ�s�,���Lh���	4�'��<�d+��U�ү��Q�r�!#�/f��.�tH����y�+��6�:/��%��O��g��-k��f�p�&�[�g�-�u��\�=g�h���.�f
[N`h��(���bN�#�d:ɟ��d�}����R0C�
��@K�ꭇ#H-DW2E$N�(�qy�4W�x����)�Vυ\Ɠ���,1��鏌f�qv}&~+�o0K���=�~���zR�gJ�����=b�,S�g��Y_��������;�j(�1�h��iQ�囷�pzS�1�1��ȞR�7բ�	��Yӓ����Vκk�C���Ǵ�1��R�U b���#d9X�3*?- E�2/�ğq
"��`�>���$|��sèJ6ȠR*�.�ki�{�01t�:�&n��-[{���U�-�8�~�%���zZF�P��T��'������^�4b��7j�"n��TP�Tc,O�IE�����|J5H�)��z�N�hy�I_R+�'�Zō8_S}��_K 1,���m2�f,�����L�
��K܁�E
�~R�:����ߙ�w����q��Xs�fK]Z9^�:3�E=8����2�C+�� ]��#m�z�Jte�?�A��^8��]���vț���ܕ��Ï���=�a���U����i����4��h������A3�l����Ii�X�Y�?)>d�y�q8+AS�nȇ`����A%;��L�������)I���?�x���ٯX��ix���}[?�6����{��?@w�,��*!*rh��ڹWO٩�>"#��
�o���<��͖D��W_�#o�W�^�����1>��:�-2a&/kZ�8����mM���F�t�]��-��~U�5��m�ޖ�q�6��*q�1�4J�辜C��5C��Kʀ�3%i�x(i�'T\���-tˠ�v*�{J�Z2��Fe��h¿9�_��6V0�q-�<��TaK��D4�K�
�̥��m!
i��{�s�b��i�u�-Doh(��IS̀�`���^>�5��,R�@�Ѣ���1�*�0'�>rql��m��MD�?-��7s����)O�PU�g4��J�D�M��vQ���������k�!��3�%x�ۯ�С6I	>_��Le����u۴4fm-/�-W'Z�t]�"���T�=0�����zJW�Z1ޕ]�<a�U����I�]j��q<ޯ�yB��t��b[�^0�(��Qq�M�<J���(�V!������q�}���OQ���-\V-<^;��M}�5��ܐ̢m��e��t@���4^g��',d�6C���}��A����DlP~��#�lw
����V��a���>�Ե��xD���T�O+Xͯ��`�_m�
0��$fk�T|o��2LI��Ꞿ��]�)�.��5 	W���-sO��k��^j��L�a��Ѓ��v��"�)Q�{��I�b��Xv"�Rٜ5���'��=�H����Vs�^�|Dr|�d�L՝��ܱ[��X��^+U6��VH*܍'���G��P�R�*���''�:BU��V�.cy��A�	��|~+ӭ��>"c�U��Jǅ~o#w����.��J��k��d)˄CW�Y��e�az��\1{"��A@�r������2=��%qg��E,��u"#)�˜b�������˧��u��-T��vZS�{���"�v�k�������d��p#�|ҳ�_�!���i�~~�h��Gb\�`���~+��ʏ���;L�H��x6��Nէ��o��9�~8���z�T`QIklB��j��a~!}x���]r��z�a!�e�
�-P��_����V"�S��"��a+M;�s�z�v}�@�I+�钝����X��:�
��H�͇� ���˨���D�=�OQ�^@������CVa���5�[u�[����>uʏx����b�-�5q�w���:`%+��V5��C�����Y{��A}��S8���	��@��ܔZ��z�����z���_�U��iJ[�f�_��������
�N[I�I���gG����\ L/8�I���0�Ú�)�&�NH�vcf@Ӗ9�#]^&f��o��/fR�$�/h���@Hz�XCZ�`v�*���O`nXr�k�%������H��}�L�XO�7������^��By�G� �:�{CKҕB6��W��1b��͊�Oc�����^�����y��7YT4�kJI��i@�!}3�$*"��-o�կ@:��h��3��g���'NO�F3�Ծ�X
�_\2��ih-ȼ������F���t���ք��BL�g�U�QMѵgH����cO�W���£�9�}�p-�����].���?"�7k�G��I=,U���oNQ|�7��oF]��C�=��ģ�n�ےV���:�p�ߒ�\�c�8|���k+n�î�1�DD��[����L��!Uu줯���y՘�b]s�땣*D
Yp��:L����\Z}ZOXb��_������ �3����` T,a�x����g��Z͇"��1_6����1?����D�qZtͺ�l���7���:)C�_͗�[t,���:dŤtx`���xf9�a�*�4='��a� D���<����z��)���2RM�@��HM�^�
G�g�T-��Z?$[2������:�-Z�ၺ6o^��Tu�4+�OC�J"���5/C��|&M���'�2 _ ���M�7BJvs{"�\Ѝ�d1�*:S-wW�����A%�F�Y۪��=��	�~�?aX*k4�z�^�[c�PqT��$�z�����=Hw���'��2�`��&Mw�$I�X�X���A�lIu�wNO�~��x�b��Xe�PB��
�q��G��H�T�h!_cm2&�H,���C���U#z�ɲ+�j��I�6;�<�ӚP5�k-E\�9�Y5�v��T*V��S{A�D7[3�O���iFTG��>��0��X�����EGu*�q��Բ��vJ�X�;�O���`^����Sr��V����6hD�$S��lV�p��f��wԳ�oc�CK���o�����1bb�(ux	���]+�-.=4�[��@fn��qO?	�H�U��س�R0���(�K�P+��~�P
����n����b�./�C��O	���ۙ�����6���J����ǆ�:H~Ǘ�H��,��ܹV�	8w�N��P�\"A��%ŧ�;(�� �Y�Q!�[m<���KS&ԫf��ǈb�j"�g���r9�_.M)�� u��`�HZ}�r�? �H;��I�@5	���+��J4�g��M�Sя�p�!g+�������DaJ"�3�'�ڬ$"��b�I"++��~o5Z����O)F���°����r5��"v
�k~�:(�Gp0����!8C�y-i���F������ɾ�^Q�	[��"�b îݷo�&uf���� 
�Gٛ�4�k�B�R=mú���h� <#M���v\[�� A7�Q����E�f��YC߸<i�Z�r�zC��)�m�f���P����O�,�x��U<��U�Ѣ��l��^x���l�qĸ�qWj �5���o���(����u�[{x�}���#+��	2u;���v��m�)8�2��-_����܁�Q�)�.���2�Z B?,�N{�7��q�/Lʫ#��#5�����!_2�=8�b�{��KX{%�zT�1�|�6.���a"��1��O��O%r��]���aj:��/XXZ�WЂвɞ���4�7|.A>P�aˑ�ֆ�?�����)Zd��ZI�&��F�Q��2Y�:�X.���%���;�<�vBWg���<	�=r'�Zʳs���䑩'C��"&��N ��E��|)��n�LX���͞�1�MǛ��w��&�x8�X�	���f�v��u�6�o\�����>/%����$��
;�i'!�`M;o��W���b���c�[���{����"x)�E ���"}�bX���bU&���7���X�V�_���I(-U\>Ɉܪ!��*�[w>X9YE�}���TZ���礣�F�Wb[p�_�����j���A����U�~�&4��r �𷬢�<B�M�=(��w��Q�
����j��ْ4��ùh_G���a;�oRt��/��2����nEڄ��vӨ$ɼ�w���O*�Dw$�`̓�V��Ũ�W��9"A{���u�J�����㓆�ޖ��H#�{�9qS%D�l�m�,}��A�U���Kwx� ��Z�n~'�9������u�dKp��rf�����L��i揕�Xa�r��U�F�����X�R���������(),���T��ථ��oW?oɇ�� �-��ѵ�a�k�zM�_/�N��j����N���V�7w�j�ԗ��}�3�Ir�I��O�Y]kDA3���툊�p�390D
��Vv�	��c��/���T*u`�������4�^Z�m<�մ��RUm�, ���b2[-��A6�b�K���M�;�n�N�mJ���(�wTHӯ�7�li�f�����u��X�,���r��w[1�Ȟ8�Q�"+���t�4
����=;G��_DO�Q���������u�0j�$\RqYJ�����O$R�a�_0 �aҗ�lz�լ���جAe��0�R�I1�;���#��bW朰��\P�����I������2;���ͤY�31�b4F+~?X1�}9�c�
�6��Mmw�2L�=�#��
�M�kbK*p;r=�ݞ5�#�=� �~���s�r"�G}�e)T/I�C���k�3�s��aAǪ�����7��a�$yb��Y���GH6?Q�B�O8��=��+[��2"�-�l��b�$���A'J7Gh|�I�Q,s���z%�\t�4-aa�9Il�뤠�����'ao�eT�I|��
,s�pU�`��)M���!x��
&��4�c����D� ���rG�zZ*�e���Er�+��%�%��o��eq���ڀj��%�m�z����,egkJP�܄l<w�������S ¾s ���-Ud��`Ӱ�&�}'Q�[��?i�}��7"�a�7��Re@y�DLㅤ�8���TI��1�sNü���rX�1��Q��{4�"�mB�-ҽB�K`����9dc}K�<ǡ�k�5��X�h=#�V??�ˤ�xʒ���XUȯGdu,~v���ͰN�������$@s��[�*�ٞ��~ݬ��ly�d��X�bAІ`�x���b���a��U	���ӷ9�	  �CTv��t��su���%��y c�c�n���g��J�d���b�oE��5���'�k��5e'JS�|�Ί%� �r�pN؄���'�������y��܃��H�ukuw�}���T���8�2@��x�J_D��Nz�9� �h,�������S&K'�xT礑�Y�7c-Ӈy�G����E�C	���.����.����NKnh�����n�5ax@g�<����B:��<� Ĭ��]�����Y��n�Ԏ5�26�����,�����XC�M\/��_~�3V�3L�����y֚vJ4X���sB"�ﯓ;�1%�]�A㎡m��J�mֱ-;�¾��-�o�w���$�z�RN]��_��z9���0��B���ё*ˤ0��S�`��z�����sN�t�R���F��GB������o?U/��r�W^�Ύ0�nU�����H����J��7�D�Kɷ
mT�r�K��ˏ+q�����|aL�s&c��9���[ǬW5L��m���X��MwmW���}ɶa3���-�ќ��*�i�#&��yLY|z4!,�5�Z�د��}��ڿql�-	�չ��Q%&��o�#,ASBQp���3*
��v���1�j��6�qD���$������/�m%m��;/�ҟIC?Ow|�5H�D�,�������$n��`��7(�^��K���.�t�i"2h�ܶ��1��'a���,e�IGv܋/����m|��o�>�[���&�e��@�n𓱺����iW�ϽG���a{o���`6A*��H7��ϝ������2lt�m����Ax�6Nנ1���>���?"�Co-�{~WJK�����1n%K4�*���
�5�<UO�u��	K0���O�J�����^pG
��}�5���#�&YZ�m~*�	l
��ޖ��K_-�}5��^�gD�d+�k��\-�B�0��L)G��9P^��/�^�x�֞<�>G��L�$!5c�%K/>�)�04���-����s������qc���,�����-kt,��p�[�<����%H+[�R4�b���;�#�T!�̕k�
�?}%���m}�ģCK��p�6�Ew��?H��a�ⱟ�|J�;<C0%��=�wQQ�DQyr�	���6E'5.`���ˮ<��jD��&T�b _�?�zW�H�Q���FK�)`�D'�����&I�����`�"����j07�,�@vp	Jbn�B۰�#W�u��(Y
��C6�Ί�^vѯꒅP��#T�F�Q��}��f:���"�˲D������۵~�Կ����=hd̗<�����E6��X3�B���$���}U�Q�BՎ���F�Gwn�Rq�c&%��-u�ܿ7�ɇl�'�݉5���z�O�(���љ�����K�S)f����h `ICW=�������������5`vO��,�"�bT>:A�:���0�A��uTLȷ��jϮM��˰!����Drl���Oewy�H��c,僎��u"4���s7~�� �_����n���ّ�?dvP`��]c��}�Jh��ՅL&�h
Rd�G)���п��os���Z�6"�se�Z)Ş�٬��F���ơ�/�9Kj�ۍQ�@%�	��I�D�^{����͹:&�� �N���y���z�T�l��������>�ōb>a�be�{�3�}�ڟH��DW�P�[�n��flm,�*=���4��S:+p���n�G֬S<�k1�Cۍ�ޡ��r˹7�`8�-7F���~��h\�8��O�^�ˀL���be�\��-�N/��7í���G;��i�;u�V���ȁ�U�f���eP)kǀ5�%�^;�͔�:Һek����|ȇ\�M��q��s��?��A5�`�K1�;�	�s�\^�	G��9��/�� ���!���\��l�U�Yާx7{+­�>�W�BJ �-���������[�6b�Lw��o^aDi�/ "k�O�ǟtT�B��V܃�j�Q��K�~�7:�����و� 4�kF���}�}�![s���_�?�aU��d	�����aUD
��a�Ŭ�̷��$l6+����xǕ͌M�Ac���q�"j�^M��(:#<1������)J2Dw=���ٕפ-Y{V�2S~D߰�=;3-5�ѱ=q���F
�$Ow���|=8"�+��q�v�u �Z���G��,��) ��P�ߤ��̝�(� �O��Μ�U�g5��>4��De��:]1��?u�t�"d�=�U�#z������������o�e�U��	�����!�`!���4��¡���ܼ�ɽ\g��8�?��R'%�ĭ4T,vf�w�I(xj���Y^��j��;�.��F��g-Ձ{UOzj�ԈaF#�;T��C��w	�*ky�5rfR�Д�+�$�����J.�Zv�>A+��]�*���6N��S�&�P�2�&\�C���_$����$�N`�r׼m��$Ԓ	�>�?~���m���7"�F��d]̔ɢS �*�)��TX�E�ǻ����`�U�_/)�n6z���
%s���I���yTb�d�$O'�eLT�y{Rp!���7*�ҋ]�S��AJH�fĩ��\)����ޡ��XP���.��� fYH@g�U���,�e%u�G͘Bw�F�f�DGg墨�k�sgG�n�ղ�{I)��R{_�hG�R�m��/�Y�=�?�WJ�i�ߵx��J����5Ր;y��z(p�Q�:���'�4΀�=O~�l?�a��o�ci��s��Ϫ���}����o�i0�q����n�^�p�����>]ajm��ԁ�\<�s���w���׳��sGF���h���yإN��U_��b؍b2�
����5D@A�N0d�*�Q-O��D��#�O�Gy?͑t}�!��P6�,�#>����P����Z+���$��t��ȽC�BGD
���G��{o
AE޸$��%�ǀ�Q0F��/�6#UCs�&�X�1o]>��٘mF�
A��XX��c9������ҳ (�!4�s��2Ե�H���J����L�!�xI�c�n����w��#U��1��6#+����#�e0�%pX	�v~)�GAt���IW��,�F1_j�����?�q���9ɾQ��pQ��X�[����k	=���	$��,�2O���"�X���@�ƅ�KĦQ9|_xG�epßr��/W�&j�}���NO:�W�h� ��K�
��2�e��ƹm���g�61�/[�U��3��/u�v���%9�0&޺�� ��^`��l4�6��1DG���b��)!��C7Y�6����D���8��]�x�DŅ��8==$$��	Z����vT�Z�#c*�*�J��S+\g���ϕ\)�hs��������8���`DԵ��p%�� ��l�W�0�Z����R�g:�O�u���"I��_����o�L�+lَ{�{������-��:�׫!-�!T����VM�-H:@:i�gkᏮ����q��ʎϻh �`�_J��9!�G�K*T��4���2�����3�=B�os�直����ж�����铆.��<!5�����,����p������������IL�����46���#
���aj��B`n�?�L�\)Of�?�D���3�x�f"Rjk��9�n�w��U9-^J��w,v�[��.��?��׊}0�ڣu��b�Y��$��N��;W`Hߗ9O�����*��D6 v��C֯11 ���ǓC�����-��o:�k�*��h� o�:�׀���ğ��*����F*~�o�G�w��[�v#��q|P��Q��gsK���m�hn��
haQ��G�c�S��#×�V��Ű/W�Qܨ�WS�5N����[H;>�Ք�'w:��B�>��B����`�B9���0� ݨ �Q���ږ|>@q�OVl��B��@$q����b;AL�����w�($��n(��h�^:[�x(M�T�x�]`֝���q�1���VαT�av˩P���Br�"�-F�Z����p�&���]����=�q�'�G(�=���L��'2[�L
ɔ�d`*�B(#Q�� �V�83vH�RZ���1�s�₉=E�w_���q$*�Ǭ�9T75��E��JyJ��Px�ϹF���׀*�D��eƅ�.��A{T'[����ѝR���"<4���)�S˺5ka��	���v#o�#��<�KY>���~�J��Z�u��;��lT!t#\���]{��V��cc.v�d/�]�ձ�7V��Q�N62���P�I�q��۞��ǹ��G��H*���2}��]LT���rXT~Y�s%��*�$�ΈXn����F�rWA�)'/C�T��g���f"�9��r)=�l�L��l�.��A����U	�>��2�w�{E;Xa���N'�5�-�&�s�+Y��� kKW�9A�[
d��i�Uy&�>��QZ����Qi��B�@��^s�w�(��n�4e��х�7�Z�ϟ������%�c��1Uwe�ub����-��?a��dHE
q��Ga/���C��C`�9����œ�����7�K�g������3�	$
|F��@`�>y;��!�k�u��h�+���oh'-8�r����0i���6&k΍T�s���%�[���8<$��~Us�pVt�/B�=�[ c$3����Jv̏���}�],��p���2�5�1�J�����0��]�Lv|�S�HE|�G}m-CTZ�mQu w4�Dȳ"���ڹ�)�2��6F�����?�&�[۰�jZ8�Z�=�ZN����4���{9�&I�B�5���b_Mi�ޣX:�Y̹��J�,�����/�B��5)JKU�hr?X��O�`!�U�ܟӪ�l�D�vк��
�`�Ц؍�N %~kt�<�a}�R����~pc��.�-(G�n�j����s�z7�@���[����j�ڒW��1V��;�,�ȡ_B��o*h��F6��,aj�4�@<�|�g���1TE���:�h��/N˫��ټtn�Gg�X�&�E���ķ��A����Ā�ME�B�{���K�.�=i�T�U�!�89#4���u�/�˙�Twi�'%D��j�G�p�t�qۯ�Sc����ޝ��������t���S�Mf�
�5P�L-aQ�#̞O"&�P�yv�X�$m�mKܗC������:8��=���w�',�����;���S?!T��v�M����
�[�mW8�$���e�����o���Yө5,�J�r$�'R="�_��ćiaT��o<���ƀl��J���.�7�Y� �%=��J�*�P�����]����ʩ[#Ӿ�BRG��?w�>�ޞu�Ͳc��@�j���D�����H]br�N���u��|U��,��lD��ڷ���p?J�~���|?֔	�V�XѨ����4[s���v�[�;�! Pl�o���Ѱ�B$�0�>���#�T��KP/�o��O�K�ҟ��NQ�?: �<�� iEPD��9)��_nRt�K��=�#P�*�T9%,��t�o�c:\�]�z�r�Z��Wg|��c�L#��أq�%1�	Vİ���Xw�O[:7�O���ߺ�2WM�@�:���þ���FP�#B�Qv%!�43�˼�c8󝝬�c��ؐ�9����~�*m�'Vak,9���f�*j�hЋ�1\ܹ�\m�x��g����'���7`��ߗ��������'=o�&��rB4͊����[]����-�z��rЪ���c,!χ@ё�0V�L�y�5��UBn9���]	c[淎��,��\�N�<g0���qaS�|�)HuJo�~^�2�k3":�O��.��j�q�8�N_[�\�mŤ`�ہt��D�9��2_,u�r8�/d���A',�96��E�"��&Qj�Ne����4^�ݤ$�U}m0z�U4��;$��9� ��2Ԑ*������ϭ%8N�{��b�[��
4��{Ӫ��P����g��Z׀�m��d�>R]��M����;n�,�l׽���V�Ef

�6BXc�
9��t��^yd�F�3�>�x�$g�t��˼�I(�y3�i��>*L����)Ґݐ6�f5��g��Q�>ԡ�⊦d�`ߩ�kg��kwD���<��홊���ψ)���Ý��4��5u8�S�nC@5?����^[�����%���>[`�i�a�q�2t�	�ڍ2�1G���{�͖ߓY$�+�U���S��2@�i���q���~3�~������	'��|�����ɤUs��@k''�m�`�����j��K��*��OY�ol�u���O����W����b��A� *����"�9�V\�m�C���b���$�E�w��?�/e9BP���D��x�*���2O�E�m+�KNH�����2�cG��ݗ��7̈́��gϕy�O��]7��K���`_�X��Ӻ�my�~�"�qSΧ�O��~Z�u�ON����Bj���K RL�5|3x����_�_�0�oɘ���u&DU��բ�ȺG��ò�o�́�f�wj�
�ۼ��E��p
oE�(0t���@�5���E���K���nY�, 0�JR���/8T7`�}��͓�?l�n�k��1�h �6�B]b�i
�ԭ���lF�1���g���(�B*/4� ��2@�de��6�G�R}���Oޔ
��;w�;��*J�c΄��4л��N��\��e���y��$�W�R�Ct8?	���6ƫ�L�-(82[t2���w);7���	L E��Dff�B�"�pC���|nkA�>����^��v�ph�p�7������jjs?�J�【�'�P=��'�U�Yv������y��r��U/Ȇ�����U��ƶ(������;��D���ű�,��.�p�w�-��������{.̗[q��Pe���jZ�,�.����H�y��ݲ��1�g{q�
�o:�
;Ma�K��pȄىd����j�4e�}g�ow�~k��%Y�E1q�$ŃP�I�?�0�O��D����V�g���tx�h�����Be"�ܫM�7h�(��+*g�I2��=(��I\�Pb����;��
4D.Q�\�cZk7��:"XBxfk7�������X�*�����s?uu���ƢO��Nr�'x�p&�`���ܖ8���iN��q���{7��͡<q���1>��F,�_A��С�h�݋S
�������P�*D>޿h�
�.?j(=�yjc(���֢A��Їy*�:O����<F\����6�K���R�*�ru�݊��"�
$����6g�S��j5~���?��dO�#���g�&3��Pi]��w����;���8X�R�q�xZLs$��䂆v�C�ľa��z������q��K��h��H*�H�� �9��U�J]J�ޝX�M$6���4ۇ��ݠ���ޝ�BxB����=������^���!�%�U}c?�g��0����1���_��ķ�U=�?+��ٴ�L�eu8??���Eс\?]�×��i�5�+u`O݁kD�S}A�حe:w7��/��C��@��@���J0L���Pa��!����mطd2R�������:�_�n}�p��Â�2��՝ꦍ6�{�1Ʋi�l���i`�xG��f��t�����E�Ēv�6ۡ*�g|㡱l'#�V	��$N�ᶫ����<��#ǦZ�m���*��Lw���t{{x��4��C[�O�^��g�"�݉��v�o�L�X>�-�:�F�8�����������+%q�6rP���W���7��7!�u�@@C�t7l؅H�.�ۋ9�M2����s��%+���yoV3��=(��]	i�P�����2s��d�{���ò`�*����Q ���3��}��(eKt��=_�-c���f1�����Yr���ȼ�| nԴ˾�T�A�̨gkµ��:@�OG���--�S�Z\?\\6t|���%4ߧ���X?i�.��&�Y�
ӛ�H���%n2(r����Vv��ݚ|(��vO95�.(%¼S�Zo�<���1�@���+���t�3O�Jw"|�Ť"�`=�S�dyy�XU�/0<D��-��o�>�����1�hi�{'����{���l!�t�Q��뭬=d��*
�_yɉ$.��e<��.2����Ynk�.�(��f�JV�{�bVF�����r�6;�7�'�\�2��*#���tk�o�ݵT9�㰔���>�â��g����/�Tpx��0�<�׽GT�״��Ke@%.r(ZpYv�M(A;Af�n3`�a��]����c�'}f�3&���U^tc�-r �;���>�
�|��@�r*..s.�֑���1˯|���y�U7��م@*��;½<(�h��n�5�&��{��~6�����N�Y���#�O�Ѯ�_X5����:��};�ȵ�?�qb�%����8Jm֚X���X���O|1��M�b�p�1|`���=��g�&�~c�:��M&!/ѼVaw͛�VBy�w�eu�︼&�E(Jt�w,�3���/��k-���aLư�8���'y�C�@;#I�oR��	�ǂ"z��-��(��EQ�	(���g�ShQ��;����#�ß�f��҆>�1<!�5K�6i��z3!	Ceժu��5p�-��v��p��}ė���jn8�y�j�<�"�+�������7�&?���9��s��,�R4�;�C9~Js�.<�!6{4�l��Wͱs�����Af\�͇���3�e�u���O���?s�$����%j/v��b������t䦨߀L!���E01��R�Ύ��â���I$�x,�h,�
��nc�3��-�®r����_�b�i�KA�p���}���?���@z�x]�=OQ�M���0�b��E��۔n�F��g�y:�b&N�Ҩ���Տb�Xh�ǁ�s���t6e��iT�Y�p���vh�l�ː��HӍC�0�v@!����E�lW+1u�(�M�m�����g��t�'u@�
1�:�Р�?O��<���(+���i�Y�h�[��\��vN��E�`6jFs#ЦF�l�2�MG6XK!l9Q��r�8LM�{}��)�AJ�ذ�;�fx�v� 놶A�*\�(��9��~q�%@�!eFG������&�'v���R*��Θ0fxW]u~w6Wo;���[�+�E1��;��"�ߝ͘�ue�>ڛNS�M���q?�������2�t�Z�]@�Ì�2�ϸ��-c^8�S�EȎ�Y;A[�C��eH�UK�6��0����_�@��<mu%ҵ��X� �s�F�P$��.����e��u�M�E��V�$^BO@�����ݪ����{5u�zjW�!�F��t���.k!g��[�;�0�D- '��Q�f�����z��RF�H�P��nz5#$�Q12�2��D[HA��)ȯ���}��#o��j�Z�T�tXT��M��I��]^\b3�AOb]�֪��̚�pig�tD�+ A|��c6]l ]e�����h��������<ӜZ�t�=�WP�m8U�dcܠ�`���1iۭ
H��o�.Wl8�花�����K�S�f=�����4��<T�ݬ��ɳ��V�����tg��R?���23�swP4M�u5'���S�쿿�s[^��D5�M��#4ҹZ�Hs��k	�����7�"��_���(�^W���|��72�Z2U�����~wD����3�H���K� J���)����m���92K�M��D�nU@�J��Z5�/���8��V}�&:�.�����)��0Ld��CuC��׮�2�ْ�[����M���D�����}�ſ,��6��A�j��>tP���a���-(M�i�����|���a�O=5�b�ߋ^&�m�uW�չX�_�Z�]�A�uUF��Aʪ�d���h��s^B�N ��j��z)J T4�fFZ���Nt=�g�\�������ʖ"]���<�$}�k����xƤ~ ��=��d�8E.���60��ȘR������,�L(�Ơ$���t����0qw0��e��5#���f�Q�����a��+�!z�I�G�I�MNz-��Th:�<1~n|}�gx�]�@i��`ǌ��L;j���wU�ԁ�UE�.~@v�S��6^S*gS]7��g���M�j2��/�\�!��YY�7�)���#T���Q�QEI��;t.?Y�_k(2���ǹ���%,}���;��xag��ɘ[Y�n�}��H�Q�0�1��?�\�a��7F��/�ς�C@�#$@��f���4�v��K����nEo�*������v��og�pY��},((�/����UEo�i���LQW���~qp�{�V����j#Q���:,ؐ�#��V�T�f#ɬ����6>���ugY@ʾ���\16P��hX7�U�r,�|�̷j�>��-�W%��6�/,}�J�|��S�ء�6��>y���{�(V7�2��Jπ���F�[5=�Ov'S���4�V�A��ƛN�V����t"�z ���:W�//;H��*���B��@�* ��N4�:������V:hg�I��\t����- X�R���3f��1J��2�듂��y���w�\��́���R����A��ByO?�vd�:���u��Qo��hx8.�%�(�]r�
��w1��g�|�L-�q��8'�+t�݌&��T�Ƙ<[SY�B=��_��{����}gi:~;����M�3��Z8Mw�7�a�A�A\����V+��[h�ud �f o{OY*`�V�~w�nb��u�v5�����t)���^��;�:z'*�o����w<E�����������׀b�x��
t�����W�RZ������Q����Sa��:ͪ|w�a��Ћ%����;��':X�f�,��o�
F���n�2$�tx�����tM��P���xeFH�n��kz�J�a�b.�f��w�`d��5\��LTօ��PA	��4�*=XI�m9o/'8��n���Fq�{�gRW����:�c��`��n����6C��d���a��H"O�U����F}wjGW���+��;�w�ŊA
���P����[���&�ʦX4�.W1����z2��>���c��-MW���	{�@���b����WX�-M���o�i��8B|���5
M�Tԋo�͂�U��^����Yp�Є�tb)rP��g(���6���յj0�2{���VFu824 ��ⷖ@q�m�t�{%Y]���k^K��X1D�ME��p�ʝ
H@��;��%~ٓ�ʘ~z�g�*=VV���XD?����P�;��w%��3F���% +���4��42#�tx~���j:����=�U��
�3ߨ�X}� UV��#� G>:8`q��3o!�*�r�6�z<�w%��G����bIԂ��	sxl�4�)�2 �������� �p�7<ݒ8���Xse�v�M �k5c�I���#�I����f�9�F|��;'iE/?�����v. ]�/�TP-�j��
\���R�;xBY�?��,\����n��T�F 2$��`�S7�O��<��^8M�%��W���ږ�F��^���b�e�ʤ����)d&v�D�Ȁc��E�w�͐�7e'��±`e�Zfwm���R> �đ��IH�K��J�H-��L��g?����ʒ�������ǖ%-x�a`2�X���ѵb�9I6��&Mmb��`ϖ������H車O;4.b�A�,�W�lS����n���Ɍ�0.��A������ͳ����L��B9r���������W��N�tֈ��Qʔ�	�R�i�
B�N�!z��C��t�z��W�a��G ��ŀ��� M`c���4g�i���H��BZf�-m2��+K��*lnmi�8��e�k��5�AX7�g�����k���l��{�.ΐ�Wj�uO� :���h�t���l@.���t�54��Pu���Yy����H�i�˄n�f�U���@����u�bD�=<OgE�A#��~���~z?��"�ؤVB5ݺ���UM�����������+�����D�J�-�ƿ������)��PId�[d�|�t$Y�ȿP�u�6�#-�%��X�nK��k�ͦ����S��Z,��C�d�*2 ��V���ГD'�`��޺I��2�2���H��wp#�t�PH�3 ��fmlZ�%\�������R~��-N p��Ŧ��	���V��Q�v�{��M����1ȂP��j:��#H;��ח���W��j�<�
+�d$���6�8=?����]_�����ߵ�~L��������Z���O�X
!�DP�L&�O\M-U��ւ�qw���@��jUgJ�  !H顒��c)�&�{�@��5`;y����#V@��KRM)�E`���su��f���Ro����Y&���iLuW�Y�N�F�{QM���H}��!�?��8�ރ���"�kwP����1#�-��u�qi��w/�cԖ7f���`�fY���s笎U���p*P�����B7�"ӱR�4K�7x-}�X�n�/�~�Qv��,c���[�%�?	�Lq'7/
�,��KU�Ro4���}hvPa�'	ٲ�ioj������ta���J�w> e�7�A�&{ݗv�"�|��/'����
ͳR�.�H/�B��̩
H���v ��[��G���z�?�4���WP�͡6�^t��O��Kn j%Q��5A	����;hԵhAeC�c��V��9ch��"?�4�x���+�̦�����̅ӄ�vԸ6(Y��O�-M���E5��&�(K@�=�h�X���I������7d��kgf�p7��wgS�)\$\{(=���^��͌^O@e��M���Iz6�fJ8tƃ��^�@��c�0�1�H�6y��}Z�Y��Z�����j5���@�԰V�ndH��)ѳ� ^Nì�Z5�	F���v������Yo:���ͭ��n����У��73޼9m0{AG��bH&���r���d�]�����)����r����o�p�h3XB�P�fC]���ln�ᒁx��+
�,��~�4��5�?�R�%�8�鞠5M��Z}��a��?/�lT�]�<}���*��K�<!���|F�p+�}��d~d�u�>�*���RZ�S&5�Ί��J�����ǝ�j�-��6�]h�Jm�Ip��(lfRj�SV��,�k�n���ZG͎f�,43U�g�]����v�,R�*���PS��T׆6QRm�f�_��sjâ��]3[,7n�M8+KW��b�x���Y��ͳ5Y��I�Y���k��X�葍�J}��XO��α��t���3M�f+9넧z�)w�9��$��.Xe��$ǱΌ{���j�ɦ�o�M����6���]����|4��h��B1��+o��Y:;rd`d�������y��B�,l���<o>�zSC��𡝸����)J+p ]
q���7�&9ۡ�d�8?�k�,R^}w`�g���f�������ʤ�<33�N�Y��i��P}�|���<��<2�4��8�"(��P��h�W�H$�qf�t!����tm�Mg&��~����j�T7L}���N�Z�"�iöƪ�^����][>�XF!h�ә	F��6��ِG��oـQ����W����yeG����HKBԠ2��L;�l�$��4�4�`�P�ݳH��Lk����7_v�����	��8�r��ZU :A�Z+=}�֒��e�-�ʲ���o���*������L��Tf�שq����3.�r��Qcq�S��
���(,��V����w8��3�G g��*%���'�B�Q����`j,������%��M�R�����x2]J6I�2_;�n�p_�r���B�l�!�����#��@֑d�]�6�@��~|�T�G)ѫ)�=�_��0PM׭r�+2�����QW}��i��@��`U���@���]�^�g�$��"-�(���T����?� �ۂ��Z�� e�o-�6���mH�����耛^l��6I�^�Բ6	�S�`��y=��t�y�ې^��i��YB0��d��'�bU�`���I�R��)���Ț^��M{ԑ{��dިQ��Li���7�:���`t��:1��h���dC�.��V�}A������q7����9�h���FI�Z�#����j����`���CX	�6�Q��l�}�	��wDi]�[��EG��HF�P��91ͳIZ� ��(<{+'��t�%����v����p���Z�Q����udJ<cB
 [���X��^%������w���)�3�Ѻh�Iֲ�����owu#�3'q&y��s��c�}��:V�"�U�=I����}]�2�bG��ߵ$���<<c٣>�芿�����Oz��<�I�����(^}�p=.{ӑ�C�둞�
���%�te2���=�w�`@�\�}gGc�w�-��l	Y�@�>dX��H� �Z#�����P���(-�g��h��:\	z���]��D_;��-#��3 �iejm��H9�L	�N��ۣ+��a��[��wWC�t"��ԫ!ai:z��MwW�`�1u��8{���w�</_.,�#��*O���z���0B  ʼ����M���te�!C��4)���fgh]��9**B�ӊ���l���@��<6�b��̐έ�.7���e�Bޓ����<�o��CӫQ�9��^�B���U-f�B�]�g������ɒ ,��ϫL���$,��	��mo[GB@BV0_��7k�t5/i�I����f�hU�&YK�Y+!�[��JI��'i�i���0�g��+��w>o44N�5�Ѣ�c�?�zÅ%R�=w\\�`==�u�[a���]���Ҭ:5�}��}�-! �U81VCL4���r�Ԇ�~�#���U�T�ؾ,_8MT����4C����(�.,�I���[��Z��׼
3��3M�+Mٙ�����+����f�����Ng�|<�8l�;Ƣ���l�M���h���氽��M�k�f)z���#O�p1���A`�c�M��<�)���Z�Cu�!�"M��M����& �`>���]�i���J�s*ڵ!�o7��
�N�����0 ���`�}�+������٥,�.Ǫ�`ji����Rs�q��zu�k�˷�Pҵ8Fb�Sgӫ0<,<3��:@�i�����A&���������L#ؐ�v���
tpr�o53�n�&YI���bSsAS1�cl&-�I�7M�pn@`�k���V�!�z\��������������{\�~�4�c�-9�]0Y�ixŁ��/��t�o�_^v���I����vQc�l��q��2ss@6`��u����Mh����fR9kvZl�E�jڏ�Y���;�����j�[�ȏ��)�u�y�$3*�"�u������T����A��w/�RW�"L���L�����w��\���0�
3���uO^����ʐ���Ҙv��T4YhQ �)�,T0��'�b�*��w�ւzFg �x�~���=I!� �95��ϐ���^�_�
ɔ���pv}HOϤ��a�笭>CMbp���"� ���z�mXu����z�٦`M�����tm/��ֹ�p���"o���6��^2_̵y��	2�7���!U�bY��C����n�<���7S�ia�R� ͤ���i��U���Kl�k��Aj�(�t��5�b��/{���>�ɳh\%�ɳ|U}�@0!��˻f�5����ߪ`�>#�t5w�?%8�����@�fO���.u��~����:��q�.yUa���#��[)ӖV�V�����X��R=h(VP���wTE�w�-������T;�WM�ѧ�q �N�}��H��͎���"�7�t�04&��8���5�>)t��"M��`��[Yӥ���B�y�L������z4�,y5�pU��ǈ`t;eZ�V��!�	H�7�-�#Z9���d3�{�"]@�#p����Y��k4�-�}7��[/O-�e���63:+"MW����t�3ڇIn��tE5	.iF&����f2�jz�(�Mma�ǤZ+����~�;KE٬�J���&겼2-ʔiIѮ��꬏�n�r#��0��B����=`��4�b�
N�}�ȯ�'2}��`V�ݘ�>d��8��HOz�E����[����#u�L�2OWʥ���KL`�����R��+���(Pqgh.:��go��iQN�Vt�����;"5�1K��e�{��Z}���T�ڤT�Y���s���!5�����V��^��m_^BMg&����"�P��� ��Y*��B��]���)��Ic���odW��p�zY�n�7��yeFG�,��t<�~����r����n��	���h�j�Qr��Y4�ΖUwgS�����Y��s���H�	�)�Z��M��d4������8��%�E��� ����[(�R��0>y�j���s�m1�+Ӑ��9ٌ�祮�D�L���:_<���?+��?�6h����x���.C*�n��f]���}7��YS��;��×�tlzU׮߆��ɱy�]����e��L
�����p���)�V��yB��	LP��L3)��x阮��n�ǳ�4:1�Y���`�d���]�oҡ�l�Ms���;�;�!���@�����}��1�}���T��ԋ����W�錴N�fU7������6i:H�MWN�� m�4&����RSk�N򜹀{g,A0�Ϥ^�I;.v�m&E��J��`��7�Q��S/p��w&�~BP$�`Q����WnE�iI���`}*������em�͖Z<A�&�C�"�CO#����ڤ�����|���+��m�MW^������ڨ����J����1��ݎ�h�`�*��m��V�ۉ�c�5�"0y7I�	��V �7v~��m);`�6W�����S�&�I_a�lU�8��*�M(e�{j�M����0YV��D�M����6��I�[����nG�Ca���euu3�HV�@�� >�w:����\x>�溭T:� Z.�d��S#��y���̓��L�é�JK����k�v���8�S}�"�}�5�rP.�n�NC�t�xݥ]�+u-�M�^ˍ��).�90"��\�L���$���������	5�|+	zn�r�^���lȿF~.C�VH�Ȓ����f�H�@��C0�U|��1e4e����;WǓ����N�ev)�羴%�o���׭�^�����).4ʂr3���i�}� Fq�w����V3��x��	�-�Y�Ԍ
O-l�MVR�A�����f|֭���3���n��b���D~�4��R�?i�ξ9�K�tYM�G<�:�;5y�of�tT���A�������U����f9��\{�S���T��O�o��B����m&��ߧ�	��>E��6 q�y��TFx�K͗5}eDs�>g�&oM�����ﮞ�Ʀ�����4M��tޭ������ݖ�|��V���a�+�Cu�ޝ$��a�㩳$�[���w�A^T��eHw�UBj#V�!Q�H%�M��t���d)��P��Ϗ�˫�jU��[�&_�����!�ת9�n�a�	�	&���i� N��5����l�1�R�%ݲ��BVqGe�C�f}���Zxr��۴U���讁սßy��껸/���<���,��D���6���k7�Xe�G==��zӹ���4��96��3sо�# �QF�VS����A�2�c�t�fR�Z���$${-)� ���3���j��!���w��2}שk�
�s�}���;�P��j:��;�t*CBc1&���M����2���w��v����Õ"2��(���L��iɽ�i	�q�1I�d��zCq����'D��î�w=��ۃ��KRxé:f�M�]��*���>���-�Z��4����

�a7`-j��֢���#;�(���JP������w�fRCA�1ESvvʫV��V�vX��,���ϻw{Q0�	/%�}��V}�S��%5��iDo�N�4�!h:���x�t���=w	ye6 �LC���v���5(�j��*�8���e�fҵ!)�}�H����k���q�{�/��0����^��<L��gWft�V�w_��RS7���I�Gm���n6��Ȩ�*���-�i�p΀�M���װ��iI=�I� 6�b�u��A^��[��dH� ����{���R����i��͚@�M5}G
o�(	�7��wy�ϵih:!4���M�u��o9�n'qA�f��bQ�3x6�*PCJ��3--:C�,w��6�52�4 N��LZ�����Ui���% ދ���=�⯯�4ͼﶚ�˩�UJO��V�]hz�W�7��2�sl��}0eg����S��9_Vа���A�R	��w�I�]��������.�wFMk�����׶Q�i���r4ݎ�{���l�Ӛ���0k�}�6��rʴ|��6א. � V*��4�K�Y��4"}76�;�yad'ϖ���o�t���^�M��c����lPb����N�0�Dq�,�nY_y�#ҏ��������%C��;��U��������1T�ɝ���j��ת�a��2�:�^1~�x�����{~�+�d�kאJ�.,�NZ�������"}����Q�޼�~�t�4�2!5u#Nz�	�<����냶zNm9�5Iѹ���g��d{MEo+qOSs���n�k{W��T2��;H��4��]�R�RSQ������9ի�4jڷ�֝����~�'����Tb̗]P?:-��+���*;M?
���Vr��CM�J%�n�./b*62�ơ8d�s�D�^�|[��߶���p�Ę�+9W���󙜍s�Ko�SЕ��R_H�O�s�X��*GJ`�Zx|s�{S>+X�sY<ܞ.}. �}��OFKy���o���Y�ih�6��J/gȈ��I�K���\>fXCU���t��n��ߤ�����5�]Ȭ���D�}��\o��p�d@4�-e4���P֍���ϧ��mQ�i��X3|/Mc9.���#Y�l�8ԫmG�9\���]���mJVe'� kGq��.d�OO���T2��H�Tf��|*�~�/�&�:'ff���Y���Jc�DeHs�O*0�D�W��;�M�\��VBPں��S��N)��T�3�j{�����}�J �Y�*��d��?Ϧ�����;�q�>��R���Hs;��,b :�.�۬J�]�=u���<�����*��?��z�3;o�+S��r���6ȫ��\�e'��{~�Y�N-Կ~VYh:�f!�U���sz�?�d�N�Z��B���9�Ͳ�K�v
��فǹ��7-�ʨ-?�a��'�C!�*6t��ӏ6U9�0��y�p��h����~��n�G{�ɦ�� ��h��B�a0g0:-d%F���"�N��ZX�#6^t�����.�T*IVa�.f��m2>;�t9��{�7�Hႚ��t*;���p.�㐁N�`�nR;	�d�7r"�y$�V]�:u�۵Tք�٬y�a��F��6qL�m6��C�<(�u��j���Փ2яw3X?{wy.. �YNM��
DȌ~�4���"\I�b,<����
l��M֧��/1�PeK��s����껖���	{�H�$� ��HQGܑY5����3���O̵��ѕ�WeF�n�71n��AH�H�$��[7R\)��?��̢���s���ä�.$J����{�d���F-�"#lذ�I6�6��t����y]\A����=R���/��g��[�s M�y;��}��Pʇ�j�Q�����^�|����ϳ%��9�n7���ln
�|��Iy+#Q����!��M$+��3��۲���
\X���.� =#������3Vp赣�8�Ϥ��B�y�n���فYl(ɻ/c6P�N��7��"��Ka�ℇ-L�wWv8Ţm#��!���}/�y�.t\��N|C)U.>�s���w��͞��b(\��M��*�(�T�dz"6m����+Hψ�x��1c����_EMk�%M���h	q�0k��e������>]��C�߫��zՀ��!{�+I�t�(F�ш�^�U��-�ze��l0�s#+�� i*fH�쐼�"�Š��:�����HIV��}|�+H����}���_e�u.��0�7ⰻ9\����_< ��}��L�?�k�PkD�c��n'\���d�[� 1)V��G?U�mJ}j�u�$l7�L�s��g��5�l���$j�)E'�����p�1��$������7]��8�S�|�﬚n�gnmK�Nx��=��U�Dj��;��+S}��m�YƶC�LR��*�z�rFl��(��c��B�l�,(�;
�g?H��M�v8vFJH[�����ǠZJ�e�S5݄��~��iO]�Ƥ��vTM�.���!�����j�~��j:���͊z�_RQ����	������F����j<6����[/a�ܓVA2��@Ȑ��;]�י=␯x�q#lT1x�~����r�����}.�5��t#�M���'=���Ψ2J���h�ۑ��&�������~7SQ�S���w-Ҷ ��i0P�ɘ;�&��5�$(��ʃ��g���22"_wGA�Y�`�~�v}��V�7���
��>W�� ,6t�^ЇgF�����@}��@!�5�bo����껥�]E�f5bl����4ZB_Q�F���F�`�ɳ�h��|/� Ez�+�\�A�mx^39kYp�h�v�, 6]�ҋ��H����#[��pUx��}�ur)G@��@�>��t�����t�Ny�=	Bh$x)����\�>�[�ó�U�ap�]����=�Lyv��Y��Qp%KS^P@Ÿ�j���uQ�IX/�����sCۭ
�A=�[E-(��My�]됬PÊ3V�X�`A:X�Ԑ�q�'W&\���/��:w;��n�5JZ�`�{�8��ùܟ}��㦊����Qv�]N���h
�N��X_	O-?߬GIW�Q�b����h�9�L��.��}�Y�E�`���}gϏ)F|>��{� π��X9��6*�8��P�1�A��OG�ӶS�=�V����v���mO�J�jՊ�Y4���w\�-�8�m�F㑚N',PTaI�ĽH;�XUtA�uӔ�>H���L����Nf�R��n
V1xݏ�0_�*a��F��C�0B��	;gt��ɩ�V����%;<kϗ ЂC��?w�������w��J�Qo8T�nW���?��+�-�D66;c�N�E�R.�l��[؂4�3U�+��i|FUmGd�3�N�McAPh��
�#4�Q�̙�	h�.;&�z���w4݊����c>�	�m�����^}V�RwM�����Q��%8�.7 �U�U��Ҁ�-�wVY�.��x��q,��Xm�&����*��u6%v�ɚފ��C���l���U����n�J�N�頦�ק�S�=���3nOＧ�B?���ك�X�*B}a�r��s#��3��.Hm]����S��v��!�hr�
ߺXwFE]�|����d�ׅtH�(�V�g��r�΀sZl���
_R�`�sr�3c0Z��8c�E�^{��gˮ�-�����wvd�t��N���']�p�ϻW�e�+�X�|�"<ҳ(���Mw4��
�o�i��(c.�ߓ��&��/����|CE��8�D�I����b-Šg������}���1X5b~5���X95�cûF��s3E��_�����L��Vo
��}�;���U�љa0T=�%��6�SY��=7*�be]d~s�IΐP�f�v����[��[y�.�#��6�:�Y�t��ZC���_�2�{^#W�քx��C�u�?��,L'�Q���i`�;��+�w� tGT��U���g}�l���h8��_���3"���hת^�!m��R��t��[躅������I?�F9��:|�X�U��3��A���+Hk�?���Ȩ�~��t�zٝ�M �i��"zx�]�w��%]�&��x�VI�nT}�L�a���Q��cq�SYwBm�Ϊ�Kj�^W�r��o�.�� M�⚧�w!��F׉0J��MwH֓���lq]A	�a^b)��+Hk�j����~�C7U�!�',�\�<��=9n��N�C�p�O�tvX��}�Ԁ=d�'��Tء��KYwj+��-
QcoO�K%.x��]�Q� d��`KV8K��Ƃ�	B�M4P�8�,�*!}���*��1�
�
 =7E�%���������;�r4�&q��k���엶g�J��E�#G�=��������JM�lbe��#�Y�]*�T�Z5��MwHr��N���84,���ܽ�!刲���y��9ZU		��n���:�g�@/n��t3��IGh����M�d�;��08��(�������k�<۬(;��^���8uc������UK��Y��<;�����QQ�u�DN��u¸�O��mZ��;?�F�>�zSQCTv�l�d�w�fp�����5riHӍ�����2�U�вÅ���+��]�3����ߟ�GL�
�?�k���@���w��w�,��^�gGW�g��k�d�>�:Kaq��N�A�QZK��6	�9� ���9��~6�K�!U�YGl<G�ir0S5�"ҺN��0��=)�᣸���tR�N_1W���FH�i���r(���s��&aﾉ<�h��2������XwHz�cM@�׽tk�ă��]�.��x��Sz�y���Vحam�*�ʥ"RX��2j�ޠ$Ǔ1%Ҁ������M�T �疋!ߌ/�D$��CD�q,�YX�:��18p�����tB�E_�tnE�n��03�9�g��Eu���}+G߭��]�����aw1�p4���o;�5n+���轿��kT��e�0S5f{r�s̪�Ļ.'�M�a�׊5��ɷN,�q,/,)��|.�y�s���J��/_:z��U������"�?��<�V��3��JwM���=v�pw��� J����n�~u��S�<�����V)��fS�J%R[yϐ$���}��Z���Y��w�>&�Q�ƂQ����f�
R�	�#M��/T�u��g}��E_}�F�95]�q}��iw��(`��a�H�����ue�KF����#97�ļ�~��}.���tJ5f��U!|�rE�k5���dX�q���[��6U��b"����!��-��M|l��Y�N׏�}�!9��	@��:DH@M����k�S5]���s��u���J�g��[�WzW8gt��T}��������$C����V�Wm:2L%�h�.1Ӥ���!ϊ��k��<;J3u���B�mݽ�Ew��F�w"�x��O�XT�J��M���۳3U�<lue]����)z$W�2�C�'m!��g]�fz5�]�����gH��Oe���Ͽ4��]b��ibq���g}���M��F}�sӡ\=�&P�H��n�F�(1fe�M�H�~M ����Q�ӝQ��n0A5KgY;$[�Vi���ft0S��;?��6	)o��xNh���X2*��#H�_|A2;�X��SC�鮈4uN���׼��ٽ��;Sk#��d�9?�*����p3<����/�!��+*�{�*�bP}��%��+u����E�6u�no=�G`�(�0��k�٠�!�A"����@W4aA�>�ڂԻ�;?<ϒ�m3)HF18]�C�C�<�h��sj�~��3z���3�Kf���3�o��\�A�c	�H�+Eժ�~��:��jǪ;�\;{�e�6����B)̞�6/bYϨ��l���Tߕ��;G�qႫ5��ì�24�=�YsRP=�H�δT.�j��ź(gy��@�p��w���rv�x����l|���g�׋��3{�s�B�hk~^�a�w��c��$��o����x�@��C��C�����r\���s��]�:�V�ي�]l������o�6z��;
���;f�>��?cxV/�F}��; �2����}vD�~���yF޽�mEGuV�Sa�wօ��t�R����D�x�j��n
�-��-�թ�J�H�]ș:ޱ�3���5!t�-F�E��Ȃ��g!:h:����0�t�2�'5�RB�(��լF�m����=�x���CC�=c��̾�>K!.T������oU�I�(Q}7��0j;�w�%�X4����E�w��v�X��CEwvy���!�H&RV����/�D�P�W]	�Q�%}��ٲ#jk�qKI{#��Я��7�l��t2�_���lTy ��1�^dAdh���^�s#��T~�=������UM�iUU��r1d��,7y��]���Q.�����p��|�w�=�ޕaG�*,��K�Pb�D���?�!=�g�^}gsq�X%��NGh�����7��Fbg�
*�"]����W������h�h�U��_������@���(u��d v��[CU:jLy�|���nV0w��Ig����e$�#��+b�M�D��n�b�Ĝ�ҍ��_�C�4S���T�_t1z�������g;���3,dA��/*q�������t�v�Q��)�����6�rd�;*��0�uG���.xA������
�����Н�H/ȠvP�l<��j:���Lĵ������!�T d�l�>C1FFU8�Нð��kr�B.��9/��!�u�������ҭ�sP�6�������b�t�)@��v�7�t�"�H��f�8I�����\HT����
�B�t'����j1,��=W��S�_P^�X�p\U�8Pd��3�*5��gd����N:$;Q�m]D{����£����3�w�@��ݿ�$/��2fR���murq��./(y������4]F�U�b5f���\PXY��ʜ��#Җ�$�r3:���'
�#�}/l�cՃ�2H��E�9I8�B[���<�{1i0�n�Q���E�t3�L�|12rmQ���nO���~�"�]eT�]����n�s��F$���PR�%D�N�RZ��)�x���Zg�{����s�b�\�_L:J�̮2[�nM}��_��m|�<���S89�T4b��h���������"ִy�Qmo�ѩ�g�䠞����h���B��U7edg<B������>��1p�[e���	��~���D@���gJ6��ڬ1������}�����Ԃ&��go%�=��g\w�x->[ /���B/�������sТ=������~Q���m�� 8��(�'rMlyS�`����iu{?�b���Fmc�3y�o
����"�X�2 ��1�<G�U�[�1N�(�Y<>;Oa��t�S��]]��7�ŗ�J�at�S@#8�����$-��I.�6�B�=kը��������SG���Q	��R���9+-�Tk�����m�l�����}{�c�����1�:��=�ևn�O��-���� �QnUy�K�!<����W�`颊f;>�O��
�h:. ',�V���Ps\=~��kQ|������2���gi}���W?'�v��{G
��+.Q'aMC�M�m&ݮ6�t'��~p��:kH����{OH����=v�R��{c�O�KYJ�Ʊ�`��_#���A����2��|＞g���
�����d�xrUC�|�=~�C;P���1q3y�j�W�M��ʖU��Er�}���R�;K!��y".H��~,ٲ�#�y�m�.���9���װ�M�ᛖ��&������ۗzkṃ�o.��R�A�u�(�g,{P�������/�J��A������D�ʶ$�E����)��^e��b�N������(Z[4�H�H����5�K�3�AS���S��'R	�e'��y qe[M����=�zqg�VM@g�I�o�)�T�N���ž:��/���wn����!�~�m�/���,���wӵz5��BA���D�z��t�������/�@��ee�֕��ΪU��
6�~��څEn�>Jyqo*%����3�}���ٙ�v�fywlg��P�� o��Fm�B��>Jgvm񦆅F3��\ ;�uRmKx>��d�87������4��%�'I�ȼ/���d�p����u�md;�V���_�s���}i
&��	�t���z�g�c�xø�&G�ZkAV�PŁ��rN{Z��1|)t��H��Ԟ�mﶋ��ٲɬN�_��}K�־r��J)h�N�!/DT��qs�	��*�g2���a4�-l=r���s�i{�aqj�������Z��㰌"��\��
'L~z��N<�(�Y��H"�Ӈ+���X�X���A�}ֹ�L#8��m���4�S&<Ԩ�/����!�P���/���Jm3�OIc����wU^��	�gds6L�ܿ���q�*?���Db�;��/����Q"$�'����}��uכ��\���U!����PSA<�!`�X�g��#	�C�)�C�>��#�=ڸ;+Z4q�u#�%�ytҗ�W��G抴i��Z#x�B�E�T*��d75Af���<@PU��¢σ;XJ#8;��aӔF�p
*%��y���[w�5ͳ��J�i�5�@�/��2��9�y�qf�9���~��^��N,Y��ƴFi�g�m2I�"�'�/i�|jZ"9��y�!�1B���
�Q������	!���CU�ՀN�U3�_blY��D=��aq�\���Y�Ux��
�붍���i��[f��u�a�:-��
#�� �p�u!���Z��Tٱ�/&�y���rA�1���Gt3�[e�R�>4����G�󡸖)�@S/��o� �c,�Ʃ�)�{��o@�OKm���F��噮ibq��<��f ����!�<uXz1�VCH?���+#��i	cG�pE��
�����nrU�ɨ�"�O�ׯ�̝�}�S���75��>xnš�.ɰ~�'m�/�]rDu����9(��Bw��%,� ˊ�6� j?�ŕ;*�\�K��BI4�8��'�0 Ԉ��I�9��G�$�&��a2����(V���4`Aq(�h�Ut|�kYSl�䮿�	;����,+9t��Q��S��Rg�Ĵ���7kh�(5�h�f���+!8��ę��n�7���g��ô��2t���uv�RZ����5{�t��Id<���U��/V�n_z��{��Ʃ���}�M��~���q}�qm.z\*�yZ����y���7Li_K[ޔXd��ų�s�$�<�J�4��u:�vcG7 P&*IX���V��<�{~�2+ē�X^Z�d�ѳȨ*h�~����[|���a�+,C�Q�,O_{�ɕI{3��������1#؟��CA�U���8R����'{-(UuL��t�~�TO���Q3�Oy��/�G��L���R�C#�c�6P� 0w��hs��FK�"�+Qy�%L}n���v�u�}�]���ZU)=��	�p��b} )�������Р2�ζ'{7	�j$���p�yߨ1�~%㙆�<ĥ����5�:d������*����n_>��X�X6L���Ch�[�Ug�-H�W�nϦ�MDg�'$[�O82Q1nE�ET�/E�G6���/F��^aIs���Ym�{y�;d�܌���s'���!�g����e�(��?�婹x�<'�6p�쎳j�k��ϰ�jPq�p\�C�ޞJ�ej�VU��
y������J�]�e}HDU��3l�}Z�̂	�H��z|<r�4;�.����w���kS��Y���a���	��(��qI�X�]�J5�l��ȑ]��f旳�֔�	H�������6����k����┅/l��6�#�Y���AJ�D������rWr"}�+!��(�'��b��up� &i���"�ؾ�[�I���{vQ �B�C�)���{C�?�I�����wuz�sa�m�����[E0+��P�����DUۼ�mZ�æ�*�˹�]��d�ս��Cv���Lx���2t�9NI���L�l��+.մ�!>?��.��h�+��L���;�W���E��Sl����4���r�wH��Q����� ^��#9�V8�#.��u�D�4�@l����7�1���\����]x�=X�)����s�|�2%�_x�qR����s�{ڽN�ɡ;~!�ed'������5s{y�;���A��@��k2��J&�P�4�у���II*D$Z!�"寗���T�R��z~��Cm�p��j>Fs=3\�L9!��u_w��4o���?��B7��C�V��/0W��_>�>�!a�WxV�|<�0�n�z�`1�0��>D�Ae�0��j��W��*�V��)۷=�aIl�0�۪Urx��[��v,���`p 0�g�J��6,u`c� NF�g�/RV�=����9��������ś��^�/v=��b�LX�B�|Ua�_���".wi��<O����'l�l�2�*Ӧ��I#�n0�=4�~��h���V����ÈP�+�!'����B6��#+��V�������5��)~zJè����8��wa��{̂�L���LЩ���|���C��P�PE{!��%�b;��qس�\G��~&�$]�+	�xc��Z�Sgі��1�h�.v�sNs�;��yA3
�r�}�vqc9��%�H!��.܎�lF޿<ތ�,��D�a�R¿�7d��҆G��K�u�h�[��Ɣ�?�wb��ڗ=��� ��N�9����'�9��c�m�\KO�#s5�P�oq.�(i�[���޸z���D�e��m�)b�}t �t41�-�<݇<�t��!��\d0#�+sj�V3}_n�����P���_ �N�Է���*N����Vˈ%��+��HXd~#1��Ϡ�%w��n^�e<9����ũ�q]oh)�40mg)?��%&��^k��1�}��� ���%�{�3\j�>n���9��u��Q��o���Ϸ,�� w7�a����'R��]�73^���#H���,ȍ)���<&�J6�E'�J�R�&g�0R�Km��L��u���U}�$p`����4�3�xJΊhnM���Q���z���2v�m-�ߦ)�ᴥ�z�A$�)y&��棏����(�Y������槂��v�� ���n����h�����ޏ�"��F^ħ�zZ_�\:��~u�~ �����Qσ`򝷖dLm��鄽��H�� �o�Kn(�m����{P�	p�s�?�9��5`y����;��U�|�F"I/��R_e� 4������J�"���\�r'|&/~��o�e�e���(Q�("SPy�z�����fuο3�6P&�D2�L�*7�.	}�{�FN3O#�f��k���o����^�R֍�[n^�(� ��.�	L|h��	REe&^홟��Q@�4\�1U���(�b�(�����פ�<m�C���h��wLgS�%KΤ�,{IϹJ($m����klֿ���f�fk]2g�E)�h[�f^#��}/�F]�`fH�'PA�rH�im'��O#s\���?�A��ti���>N����&⺁�����ט\��p�b�C�i�zg9�;.��P��a��Ҭ4��JP=��}yʵ9̔�� �!�"U4k��t�̆kD���+��U��c��9�����]��3�n�E�w�J�HP7�������`|U�m��J3?"�)5�����ڼ�8�ɴ�8����~ {� i}�IҬ��]'a�?��R �_�8j�Z�h�(���2�����i�a�P?"x�a��%����F~*���V�0��3}��y2��g����%B�ىc�ݸ�a�B�!��-U�G��սB|~���m#7(�9������=���:W[%��8X������qc���S�(��ͻ/��Q8�>��p6�D&� k��Am�R���
k�7T�NX��~�S�ݜkȬ��?����G��I�2	�`��HI���,� 2-U��(n��qnx�����V�WK/ґ
�_ȭe;�_[ƛ�ʨ�JAAfU�������:��$�uZ�i`��Rf�N�>�9�w����E-�,��Y���2U�ߧ��(��\_���k���63�qv.�/���J!���	=d���2 �yy�w1J]���~�q�e:pv�[��B%� ��{����U�R��E/�X�P,��\f�k-7�Pgzi�'���tQ�·n��#�]����0
�R�Z]@ITvH�4���{�D�|��!.Cp��*��'opi!h}��:xwdP�]bi���c�g�Pn��Pڃ����0rQ�<��Y`_�sGs�̩��y�B)a�U��}�i,���i�&�]f�y!k#|�v�I1���Ǽn�9Q#ڠ DԂ��T�:�rSB�dF�qN�������(�8�Z�w�ڿ�P2eğw=?�o��G��������bEG)�6'� Ҹ��EE��������ȭ�R�0�L�~!qp'�fcl�>�9ef���|� aM�v
�F9��w����ˌm�?z}�QH����h�k�qډ��<�������;��r�E�L�P35͙��J���D�T����f�nn����EQ��9�+~+f��P~����e�[&*���5��n�9
h�xb�%�h�&h��(W$���o�v�L��2�!���2�[j����O�T���Wd��G�x��U��|ܹ�s{�&�v��:��2�#�lp����j�E����d�,��%�C-�Q �VH1V9m�Z���\�~n\'�_~!ۖ��b�^�"]�Sf�j���M3�)PG�ApU)C����$�&R&4�Aiu�R�⇍%�2��t*q�H��i��O����^F�f�Е��N���.��k҆#J>�����Q#f�M�X�J������U!2��W��7A��z.<�Fk��}6��5�)
�}�<tL6!���:�A]�,�3�&K���G�b�����,`��)E9�`�m�����/7�*B��K3��O������v�K��
fI� /99��랏S����3�����%_��wn��a�)��ݪD�Z�YE��� (���T���"�P��Y)�o�ø��~
U�J�2E�
��9��V��Z��Ez�ܼ���`��n�u��j;$-}�
$�y8���Ů�[�rX���{�⩲3h��,�3���	��g�2M�B���b 03t�[��֘����v�e�l@P�)�W&���ٳg�O�D�+)�����8�p�~Zu�s����B^�\	n*�3�,Gy?��gH/&��k���,���x��Э�W4Q_�-#��k��R3��?׀Ѱ�5��=�0h�ov~?E���V�Q��+d���M��9r���>����ؙB�Un���b��s��ݦ#7�A��,�EWNx绖��X7fsdR"��'U�@]�	���Q��o[#HJ��N��y��ǉ>_/�\��u��<ܳ��G^ � ؖSlJ�Xx�W(d���3��(�2�HO�g��qj@��Kl:2BMĴ0�ŉ�I��瀳Uk�W��)}�������>D�~`�Xj�0I>`��	!.�<ƃ���=sH�=ֺ�F,�[�W�+X�my�y�N�_��)#�u�g���d��j�0�t���?���~�:�z�f�3�pb9�x�L'���}�''�o�ecf�yQ'�%�Z��-o���C��B��i������\qEr�!��SQ��K��ŖD�7c�'�d �_��T�V��ݨ�Ů��@�pԀ�'U�����J�����93�A�4ȷ�l��9��J��z�n�oz��%��vsrr^�Jk�72��jb��0�L���z���Ӭ�&�J֔{�P`�F[Q�'�(aW-LN~�S������Wkews�؜�b�Rf^"ѳL9:��b9;�Y���#q� �a��9f||E���k�n9�G�:�A^��u��Hߏ��B���/7t�y,���#�����]�e�2�?s�Q�z��	�xvA*��)��v����Qی�=ö�-,D���S��ɶɁ��uDUE���<��E����=���S�	��	����DM��)�Gk��9z^.��j�t}�u���I_-мk}RO�9��9�����i��;��j8���~�>E�S�m���(�����[j���83Hy�Ro6��i�[/��it�2*o�����0o�W��i�=,�$�c26ۤ�����jM�$Tv�H|�:�z��-/�] �O�/q4V�c0R���)d6|.0����n�L=���<u�9�$�f�2 M����{k`�.�e��^1�@_�F���k�˗5��
/�����M�����~D@,.��ksL�w���ߩ�m��T$�ݟY<�Kl������~���fs̆�^��|8��Y1�v�W��T�tMg3�ʜ��#��������̓��Scޟ��)��FrN��R��rΌNj�Ƃ����Gsu�{s��
T̋�����Xѩ�����g`��a���0Ƈé�[y+��[~��7�ZPt4�<Q�E�j;wa����e�#�f'��'m�>�d
ӄ�ޘX]�ԣ�<��Xni⑖F�J������y���>�xB�.CTF���y�n�Fٮʦk��j)�;�i1����N�Nv��QJ����w�h�v���0$��OH���61/�����BǔV������P��s}���On�N�������&���x�/����m-$�)Ն �V��nw���>bF�5=��4!R�l�|w&����}_����\�ZN��7�	,M�u�rU��$���1�2(QF��S�Kjۺ�A��+�/4jV�������k5(]u�[���4Յ�Fd���z��wX{e��o]	�#ɟĥ��C�ΰ�o}?g���K�$����2v��M�\OU��EШ��/
��.�^90���	'�Ȭ����p����R�x0�#��L�+���n��\������sQ1"e��5IL�Y���W#��z��Ic��(^&�w���y��z���ţ���ϢG�á��C��d��5�G������|@tZ�f	J�8nrtzY����N�Q��#�w�Y͠;J
;�:��o����!��Ui��5|Y7�+�??�_hVQ��_���O1tkx�b������Oj�I��k<4Û�6�%��.:]�Y�2��8G��0agX���Eг���j[5+����͢zQ���I䶋F쮽��D`3,-6g�i俾DL���@�8���f��w�B� ۟��XUeԠ� d�N�=R���n�B�+C�����ʃ�]��٦)��4�2}�>>�d��Fj-������o��^"�s?|�)�`�<y���s
�����Dޫ��ބ��[�����m�?�U�a�D��j맛Y
��͜�r��!�F%�/+3Е�쪂���pE=�y���L�Zv��B�������oq�ꅣ�_�^�S֣>C^e�xV�вÄ1���0���ؒ��݋ )M���~�ͫ7��b��N�'9�׷����f~��W���'ӛ��U���.-*f%��ӕ�k���#n_�j+�מE��9�.�S�D�Ha��H���V�!)HH���`b[���� |CUd������rTy��i�ٍ,��"3FI�.�ӄQ>,'݇ƾ(vr�� ����%�0�����xY�5F@dB��v^�)=-7�����[�B���B5�����~�c�#�Oμ���Wr2.�Z����^�_ B�6�4����l�K�'~�C��:[P%�Ů���5Q�[�4ܟ��5]�({����N�w�*���f��<D�2����aT?�[r
�b'��F�Jb��E�Q�E��� ]oIf1������o��foؽ��>��,��G�S-s���)��b�Je�n�d�9�T�����Y���G=W�"�f�����^�G~
�8�6��x`H0G��Wb�L`:��3�r�EJ����).�T;�����cp@Rȓ�[��F�����������R�A���0��7V�|-�u�Ozi���#� >p��P#v���r���B*S��S;� �c(������iQ�U���Vs����a*��rM3[�hX��j~/\q��P)l�Zda���}͎��<�S�rs�F�n� ǝƳ^4�����z
Rb�ή��wd�IF�~�=.ĢI�q���g]�i�J!O�J�$N�?"o�9�?^���p(�H���栉lj��5��$�dj���f뼱���UJ��[��H\j� ���AY |�i�}|߲^F�E)���.i`��7�.�sj��z`����A^��Uq�����'��GC�_XH�Bv�Lyk����^vܭJdE��(�������B��#6���B|v2���&�����Z!��&�A`X̂�0E���B�
�>&{jKC�#p�.�8�V��L�e�4��;��Dݑr�Q���}��.�J�h&�(n$(x+J�D~�V
}�a�h��[��zA�&!8ڇem-�z�w����������x] ���z�3�0�2	@��6�9s}R�jL�Iۿ��.@�[E7�"�X�GR��#6�X�
����sP�y-�N/�Z��c���<��Q7�{[> _
�Fc+L�r����S��
-0[/~�v�L�>x���P���{��,=�i��8�e�/���=�Y���!�`�
�g�͛�U�9$�ۼ�-���R�@��������I�K�����mGM�,Z����=.��{
�͂uK�Q�E�jݥ5�u�c��c�r���|�����r|}�SV%�j>�:v���h���ՅR�[oA�u�Ҭ����C�G�=��׵tپ��2�8"(���I];�=K/d�_l���		p¶n�ѐ�V��g��O,=�5�g(�x�y|08� W�n�1�]��������>"�k&+�����K�W�����>!
�y�d��]d�֚1~����w�ğF5����P�0���+��N�#i�
��ȹ�̔e���n�1�
Ԅ|���6e*Z �X�qr��x�}ud�cB7mp�]�%v( ��>nRE��k��~l�y2m�f���U������}�M���Z��Tڗ��+�����U�����BsЬ�8��]p���_*�/��<Z�0�}��*4����FH�"�d�
��@�Y�r�p��P��'T5�k�ƍ}1���*�k�p�����ex�ec�V����C�w?������̊�ٍ�3��S�н�o�8ֵ☱��\�h&$*n���)klx�Ι��(GO�P;�=��Փs^��r���+ya`�����"�e,���ׂ���������(@We��m%`�P��	�]��ih\��$5)�ux����KD"'h��La��$xj�%�ڕ�����I̩J�Z7�G֏=���O8)���+Q=/"�D�ڍ?i����B2��+�����tQ!�nY&y�"���[��׫wC�!j`��h(��
��x�a_��t*�O�'1���!�{��JY��B�\ W<�ͽO����@8�zct��;�C��y�6'�}���+��c�LRSuZ�-�������-*�X=�K�IYY���_���2O�N�i�:�]^$'\�<�/�|\mu(����	�S�Ǎ΋��I�\����>qK�#��p����a�e�ct���}��H��C]�b}?ZzN,��u7\福���j�È� � �C�O������+���1Czo���hg{�I&�)V�:�_?0��J�ʠE�?��4n�r�?~�Q�a�I�>f�L]�E��'P!���66ƶ#E-�O���=�K�����U���Mǯ!������IF�q�(��\ޙ���;����K
����ԅ��u�p�6J���P�����	���V{�_���;Ԧ�t�ޞ����e�z�CG�;Q�R�#N����uc]x���p�s����|Wq�)���kJX�ȔR�IN<���M�[�+Q�#e�w_9��4���m3Qv�[$"�'g�7T.�P�8G�r��YS��z��(a�	"0���ӣ��cL*���0t�2�Qͮ�~�ƻ��Fy	��S��1JB�Ă
:���D�iU?�]�/���=Dm�#cB@8PR�P�&�;C��_�:Q��D�c'H#�IlYA�P ����1���k�15�N���sD5����lɲttm�N���ِ`.,���-$�_�9kW`�T#��p��ͮD�Mh��yW{��V&����y�U�~ W�\놼t5!��"Z$D�mt���?C�4UC�1��y�>��Q�k-��g��z%���J='޷��{R�^��nN�V�7����5;U[�3=��T�a�D�|���� m_nn�Tr9k�[h�'c������A���_D��ЈOM�?}�O��t~;��8��:��=r[���������@c�C��q���γ_b>�`Xw�N�U�c*%�Ț�`�"C7Q�	Ē%�֙CR���*e��QL$V��4������0p��-�=m�u	=�ҡ~e���������yhx��_�^�:0t/`���g�k����j�̂�	[�nTg�������hu��W�[1�noQ�B?�j�#@��Xp}�)�#j�T?�S�p������5���e��5�E���+m������ƫ B��W8�K4c�$5R**
$q �VzY��*�Q��EG�#�v��e���U��ӷ��"5c�;^[�o��;�m�#b:��B��'h-p�La�aN�Y�U2�e�	v�{P��N�7k$zT�mQ� ���Մ��&j2͵��o�HH��H߯j�0VE�.������r�VI��d�;���^�1)@^�Ρt����^�o#P�
^�fcF~.��T����9y�&`j���h����._��یpMCU��,MJW�C��
���e�c���=�J���3���,!CR@��?�I�h�Z��[��������ZX�/�G�=]������J���,��R���b9_��y�P�py�N��qvD�}����+���"�å~d��SQ����u�up����v�:�ֲ�p*�%pH#���|�����]z2��9��I��,�I��$��g�m)"�H]yJvX'W����X �-�����쓍i��*���3}����٩q�ٸ��?m���w�����n�W� Z`��Y��?N�!|�1�P�xK.�i 	��5.-y�?�\J��	�?�+�����Y6۩��M�&����C�=%���Nı��P��;:�9�"��n��ѡAg�o�
]d������r�
V���C��+ӌk�浏���D����,E.�������aT���m�m�3��`3ϳQ���mjr�qĒ
;���aH�W�cw�t�#`��y>�B��,�C���d* �c��'��r���߆�D�F^��A(�cC�cȳ[�=��wՏ���^_?��m�� V~;�F�|���TR�%�m߁|�6$މـQ�:DArd��l[�����ע>7�\E�VP�P,�~�@�[�T�B$��U����o�B)��V� �$k��8=�˲����������}��i���v��� SI��a�!�N?����Q�� ��P��\�ĕ��{Y�)5p� ��p�5�A����m��L��j��[�,��##�vd_���bI��2�O�l�1*vDH��h��O&:[�;��⑗Ó	|�5�&�s\������x�s�$TW&� ��'�Dm�m>���K��x���*߸�����
4��{j��U��ƿǃ�
��Ԁ��,,Q�k���۹�n��GQa�)�}��76����|*�G�?'��o�����7�x���-���U����gI徟U>�<i�/�����jÍ��T��`AU��]��
�hSG�e��y� $��bojE ��T�ȳ����~Oe괙���Y��O�F�+����xǹ^��թ�$eU�r��i�"O����aRT���"�2��@&���^RP�����X��)U�/|Kn�lTZ� ��{c�#��?�I����B�ڌ�{�,�Gj$���-���_f= �I"�'��x��?ꛆz\�����Om�Q/��awQ��M��b��2A#"n�(�l�2���,������X�ԀX�V�5"��Y#
,_���� (��#���H��|�Y�{���QZ9�?J���!��P�Җ�.��8x�C����ȸ�.��B�����.��6��s�F���4!�΢���R2�;�2y�����Zu�J�g���f���`�w��Z�bڄ�`1`Q]4�@�d��诨c�}E�뛋l�㍀2�r����&��&�ioꠟu�$/�ÛJ��V��O�'�G%]�g��ے�˱�n���L�ȓ�41�n	�lk�P�R�6��B پ׷q��*��"ͦ����k�=�R��~��4ԗ�Z�F%����5Xά�V�~��n;E�����Vq^���P*�T����q}|Æ裦 !��Q�z�L5�"Z�l��gfu���,a�[!&fq��$Q�O�C��i�M�,T�,V���jc�\�J\ܞ	�E� -�V���ըn#�p�d��|��>>׉��&��|�VTIg�IJ���x��%�6<�X9s�̶C�8�,����>�eI���r:�g���G�S�0!�Y�R�ݜ�;��8U;Swu�Å"J��@�!�������Q��z?�EU����V�zCw�8��D��Ap)���h �Mlq?Y��U��/�~ߡ���/��:��~��OCS�A8����2�Q�u�R)�O�I�4�'��e\���֡��E>���+�=�:%��EZ�+�b���q�<x[q�W�H��X:�'�E��>(�˅U��G$��w��(����'ZN��x?d�	���(wvr�
!��B%��Sg�Q�L��V+O��<�m ���!�H]M�ˆ��b�qY�I���(�
���A�M�����r}���t���"	���b�@tki$9�][�O5>,�b�[�b$ਔ����`Ԝ����b8S�����+��^�Y�C��ДQ����3�Yhvy&,�!=LWQ"/�9��V����Alƫ5 �դ�OM{	��Յ�O��)~R��B�Q�e�k��q�R����pC��vi��Bx�K<B9��e���boC��p޾��W ��G3$6��<��{y�D�k�9����\#*Vmx����m@��S%�ފ+���2��^����W쩒1�O⺀v���u�L�Hr&��i Q�+>l�V���<�L�Mn���mp�ϯ[���I"}��ϼ������]��Y$���7��n������>57�a-�+����q1�g�U5�6�{)Uq�@�4����Y�}ϴ�}8վ�xc��:���۞����x,�D�y�=�.�k��*#�O�O>Gs%o�M]®Vj�"u�,�.�S�23,���nw����b�Vi�<e�'�i�Q�k��gqb�Q����u��{�����c �_��K�\�Y�x`�_�5j�D����`Kio8X�=q<׺T��n��a��|�<F>��3����r��ȋ��tg#ˢ�7l�:�M�5��,#�2�q�Nf���4K��=��]�L�4�H8$
.iiJ�%a���'��cY�LZ(�t���s��=8�+�u������rϸ��/v�gA��gS���	�p+��)7^���	J3ˬ�EԔ�P�6 �$��bK_�{S1F`������`2����\Ǉ
PÓ��2����)�`A��m�*�X��0�w�o��\`�ԍ��EJJu��槓���u)�J���w�0|���TY�=Uӌ�c���3)qip5w�66̸a�?~�� �A�����*�yyf���?�ׯg@�E&�"t�ݽ^wh�d[V����՛�����7��N�7�B�g��w�$�.8���t�L@�Wun��ܤ7����Tn"z���WF(��}ޝ��[�����Ww�JCD��Ǵ���X1�W�����3��e�
�R����8������'�>�CR̐$P=ٷ,�p��}!'������Ƒ�v.U��};�7��E6��ɛ%'<s��kOJ��󺜺:#BY��|:h(�x��8��ϟ��y��"l/��F.n��+O�Yxw�3�U]y����ig�Yv��OM%f�TBx"��j�y\u���#\,<!R��Oj�M�o)ˏiK4�2(�۸���v�]��4f�׏)��/�I�5��X�����~��M.K��#/�f�x����h�z��J�V�JpMGC21D*�!�ߛ�T�c��Ov�n��k�)�?k���4���ɲ��m\�61h$�"�� S��@񘧀g�x���}8�&��$���E�dj��J[f�����M�2��n��Ʒ�;�U�/�U>8� ŭ�䅩 (��?b}SGQ�,���I�P�9��^��MC�xpȪ˪���VT��C�<�m��xM&U�!���ɸ���s�b����U.�8���1���V���X4b��;Y��4H-��^g�<ݷ�ue��kR��XX��ɺ����;I㷽�YE�NJf)��6"�m�迯���{j���������X���OB����t���������>l�I�����'=�BbQLR
I,��A-�Y�,�S�e��DO�����;������$�T+QV�/��6U�&Ȯm��Q�F����2�?�%g�;-�֒d2������#V�ꆣ�"�	�.^��`�O»	�KJ�<�z��#m6u;�߀�Y��^���L�Hf�Z[sQCs���Y9��QX�x�h�Fn*fA}��K�r��b������J�<�ҟ�.|R|<�	�oj��y����������Mt�s$�-2w� igXOH%�B�F�P��%:b�֊+ ��,�2{p����� .�T����@+t��gbՔ>��6���:�zѷ�Jm���o�)ŷJ?�O ƿ�����y�3��n%+�s�Q�,1�D�Y����R��j-�(A$� ���f���D)��Hk�(b�s�`z����!������5�%�rLT̀(}ڜ��F��_ݹ^w��zۡ���1|���V7�*'���h��F=+���ת%/�	zk4��Z��W.E�������F����U�����	������)�!u;gP���)�VZS_J�+�~����U��Nj�S��D�ORӤ��܏������Bq`"JC�oJQJTL�1��8��clc2d�Z)�6�)��'-24���\��5��6������J�y��Oʺ>����_mX6a>�����ȓ���W��2W�;���M�Ov{����$�'A/��	��vs��Y��YA�Ȟ���]��L�a���Hȼ�ly��dT���N�˸w�Ŷ
+J�a�{q�"\/����-%�.��%��Y�]N�(���qiN�=����������~�9���|>���<�<�
5�����6S��
��mi6Z�1U�^j�&8����p�$[V��<��/�\:�2�l8�@h���a\��O�o��d2��@T(˖�* ULbϥJa�yгXС���f��hz[eӶ�?c~���29o`JV���b�$���j���Q�u����
[����6S�0.��g�=�X�ٚ���f-C�{�t�v1��LKx��}�����~ ��'�5��pt�
�BVR[�$����3z�o���tp�A�{S�@-|�g�ȧ{��|jD���Z�J�s�Ǔ+RQ�,X���Dm�_L�Agh~����l�9@���&Llvd_�YUB$N�WJ C�ɹ��(�]�͋�m?�_�����!p��V������E���/�.3-]W�D|3pl~�����ǂ
&��$X��κ�󥛏�0�2E��[�Y]v�I�u8Iz=;��1�K��қBB������<���~4��x�AC@!������B	�T�\t��ꟕ��<fGQ��gS5�p^�j7�@�%J�@V��T��}�_��抸�.�+X(�~D�mE|vm)�
���!ܮѾ7�:���i��yՋ�	S�b��^!D������B���y*ǰ��c�,����Z U�\�\:~���/b�=c�w�s���o�-�.{����+�!�Y�B���qٽ�a-��u�1ul�Θ�p��NΤ�kS�?.�c����&-�GЄ��T7���RF�������K�2k{?d���r���lAom^pn�d{f'e !����;��BaW��q/��Q͒Q#yb	�*��$S����A��'��D=;��6�G���&�m��Ą��W$|ͨ�81�n'�/7�
�Z���O=d�y�l����ؘ�����6bX'O�����=�@���D���k"�E	��6�E��3� ֧�;������c,zvֱ����n/Y���A+ː����Ӝ��'S��l���=׊�,����vN��\�a7����B2���e�_o?��~;��_Y<��li�ws�������8v�/|[,�72i��MQ�EO���p�N�;�3|����8�E���GCHvP��08%��V�^�i�qtfJt�~g�ߌ�]�&+��Z�o,*ԟUn�>���~����h8Rq�řJ�������pY�ă� ��bV�!
�"�L�vut�-OL�A1 4��T����������NSL�D����/Z*k5q!n�㑘R&fXZ��l�ޢC֢�rq�n��+�z���:F(���ωd��>��\3��e��ʜ�ɰ�7��jb�����C%'�����[�#zPiڗ��@��,�ABݕ�0���ۏ�^4�g�OQ�'A-z�	>$	<^�/PK   ���X~�`
C�  ��  /   images/4249a833-ad2b-4779-932d-e559dc915ce0.png��eT�M�.�n��]���=�������N XpwK��	�.�;��}���{��Ͽ3�z�=}wuu]]U}���TW��D'E����T��ք��/���W(�iYn88�j{))u))juW{'k88���o��ɋx�'�%�i��)����p�>��|n�M���y�`!E���Q��� A'*�ފ�+-�L��+������v*�P0p���5��t;W���=��.��<��$�Z&��ʣDFVfƍ�[��4"��	�^z�O�H�	�J`�������]��8f�u}aA����q�2p�:_������(�!�>�}ߴ�u�niK�s��iC[� �ӷ�u�z��ېQ�2RʂƉf-�$HIQ�ۜ������+��%��T ��B��9b#1k�^�L����F�I��0p�v�$���WS�L�����"���ėE}��i�"��9Η<����L��]�O}�;�B�����Kw�Z~����t�8�ze����SO�t�BZ8 �����;�t�6}<��\��܉1?�;�q63�k���J�5�\V����S�l6�n{
��1 ��?fss�Jl��m��x|q�qA��ᏰC\�
���A���C���
�P|�lVU�|�A���+˱��+��@��Р�a����a����%�R1�O�s��-έ�ʌ�=�OCtbSO"z��YM*-�gJH���A��Ȳ]ecXB���T8p$	��~R�\�Gӣ[V.��5%Hj���w��$�x���O4�J(F�9/&�/��\:�9��yO�8�P:�#5� 6zx�bfJ�x�o��%��I���$�K��)M~*%k���P0i����M�'s���¦��܎1�F.D���'���	�[��a�C`&I�U$��/H/���g�b���"�WTO-���������aw��,v�KG�W�y�v�/�/t�HZI�_A��hJ���N�A�O1,���<<��x���$�"Ũ|1����u��~��o�3��������-���ɱJ����m"��D��k�` p��1�_�u;�WAsn��qr#���7��N�r7��ΐ��t4�]tV����8B�B�{�5������#�"��>[���f����ń('�H؄(���e8����G���%7f��8�Q04%'�&Y!֓���%�*[Mc���& �h��H��o����5��� (�npo�gKw��`�`vRõb�+�D��`M2׷�l����گ��5��+܌ͥqK�~��j��V�����L'��/��V%)�(�~+�h(-�z���º��f͒ʖ�G�.�B�ܐ����}���.a	o	Н�|���=]ݠt��G�E�^}O�RQ�R]E\�Tx��Ye�OT�lx�ðm�"l6L���ׯ��|�������5-��ߡ�(�ի$UX��Y?��b�"8&=���_��ِ��
l���d2�Ð�*�;�mqU�Q�T���t�,�,��Ќ��o��l����������������j�%L�'s'�����_��&��-J-ߎ�T��[I��P�+�o��(&c"��9#d.|�OO�\�S9RF.FUn{cN����㬭,�e������l��;��&�-B�O��)�;鍴D�/�F����-��X[ZmU��M\�N��ᮞ�Ő4�׶�汫����U�Y�	�/�@�lE�B�"S�.��"� ����8O�i�f�����j�*��7�7m�?��BzB�?'?Z|��E�6����n����O��(��ƹm�y�xLڌ~F�'~�qSd8fT��D�_�:g>��(�$91�y�m}�4P1G�yt�1�_ս]�`)~%���I���Ͻ˸�|4|0�z6~�O��"�tF��?4��G�D�A@�AAFIE{݌1�y�*/���g��U��<]#����#����ʍ4[�������`���Fp��G/����Skʑ+v2��v3��^B��m�����_:Y:%�<�<M<�B�Y��>�"���߆�#�!�ͣ�س�����q�~w���Ӷ9����x&h���ݙ�'}R��
�
r��ItId�P۰���T���Y�ĲR	����f&g�C6�$��y����%}�g�V�3���й�z��P��E�E�����F���b=�����Rԧ�օO���wj�Vך�>ӹ[N����E���F-�&�$v��Ԝ�[��Cff����|�X����ct�|�;�֮a���ya�8��b`~4w0Zi�>�^�>�:�9��6���	���}{� 7��� 'M;�#U��:�:�:����_\-\��U��t��w�=q�3aA�V��z�>%��K�<,���L�۫x�	�Cʡ�q�����5D4��4֧����������ք��u�P�R�VV�ة�0ëʫ�߼��YM1-�N����y���Wٜn6,�'e��|n�g��(Zk$�t4��g�����E��\8\[�����:�w��Ey�:��\r&  î�^��}SE��[����}ܺy� �+��e	�t�x$z^qTc�z�J�q ���)\��T8��������������'�_ �c�S���5DtП�֭�n����Y�RN�������p�������5*,������o��[�M9�1��Yd��������%נ?��X>;̗<{�7x�{8��ތ�.W�hC(��� gQ�����d�0*�����7䧷�[�\?��Lc;�����X��p=md�	��>�ù�#H�!z��m�/f|����χ�?1�@�:ՅC Ù5�׋[�yf6���/,�{���V�s���s����y�r`�� e�s�9�8A�,����Y�uI���!��FY�+ب����گ���I�a-xX�'���,<3��pp�pH������I���?OĤp8TXV}~ �w4|���i���IjI)(��Z���.�v�^̊��47yO88"��
��I��������WQ�tu�4�r����qv��~QaX���˜�����S�G��?#�a�n.Z���r��WQ��r���~����M+�NMM-�ae#�)-��8������0  ��q�z�r�{��������6������܇�œ�I�;�������������ws�O^b�������"k������_�`r����������_��V���v2��w�a�!���V������*��Jr�����ߒ:��R�ΰ�^��{���?_�������/���\��g����X�m$��Vӆ=�u�9Xe��	���D�^��CNAZR���c'��w�ef�Y�5";��f!�������y�Xq)��-2���=<4�T�Z-v/�8�휘��7��%mk�,Q\������ �"�5]^y�㠋s�Jq�U´�<�?�9%I�UZ�0��=�(,��#���������p�{`����
��Ћ3����vHjq���V(��S��
�M�����')!])o 0����v���!�X��Q�w`7�n^����]���=����R�aZ˟�|F�A�ޤ�`�o!&��ė3w��Bk�5��_��0#�JŴ���ǔR} L̅8��ڹ
����(:{�n������G�������֛`�{��[���t z$\ć�gF�]��آ�ל�>Y\$��y܋(��>y�C�{�B,�{�e,�"b�G`Hĸ	�pS]�� b�������	�n>h����^�	�d^�)�q:�����$O<���r4�-2U�a�Sq�ڸ�[�����&���ʌ�BT�9W*�p�\�pWJ�PII "���W�8�EfW�gI�{�gC�gl4{��Q
�O��m"x�%����q���g�b?}[k�"���LBY�S�䋺���>�ͷH���O�"�{�G����Mm	R�_�~7}���¼� !��$r��H�D�����`e��5�*c�p�f��I�z=��CU�<� 0�1?��X�vǏ���/-�ډ;�bu|J�&��z��_��-7%O˵q^+_��tW��<����$?���u��A��s�M�}�Ӷ�ߣ���'��/V���K��ػ�7�K^����;�e������G4u��}6z�{^��6׈U'��z�B��?.�����F�;II�)�($����?=�	ؓ{g�3{�~���!&e"������3��B`����˻�>�����6#����C� ���x��pQ���J�
�0 �`kP���PDaTڨ\�܇iY>г�0鯌�Z�e�%��H`;�%Ks�0���T��Gd��54!�r��ݐ;o8�F�F�צݚ�-'+|]t5	�hJM'�Z %����yxD�(k'��O���*s ���=���3�����i��q�d�1���)`�F'�
�	�+S�k@�%�҂N���d�:
��9�N����I�/Χ�z����r�\��ą
��ŋ��#W0�i�0�h+^2����2��%b�)4�g~FIFu�Q�ڪ�*ZzN��E�ǟ��R�����n~�'�'D��`!�_4��?q��Ĺ����x
���:���ǻ�)O�o��pe/,��aZ"�%�a��sn
�DN�"A��CxN�	D�����bU�.ꃂ'�M6k��u��O��8&lm���Hz�H�/�v��S>7�c����k���2������u�MC
E�!aPm6�թ��{Y2�~��A�4!�폏�m2��� �ϕ=�F�O�w�E&�rp8��NrFcB��s�Q�2%}U�Y�Im�0_-/͹���LRN2�yɸ
�:9��r���'K���*��9/��$��m�}�j/�
�$^�^_����H�%(8���m�6��X�o�
��A=�P��,����"6J�נRRj�TW�] + 
j����zK��<U��i�)�=�6Ž�i4���r�R-5��1ٯۿ̻�|4�K���|��}k�4�͊a��F���t�x�	�?�U�>`&�$��DwD�K���^&�׆v�ѝj��Jݙw����t�$Y�a�|"��f2��A6�X�%�]�\^��]���|)_�V���縠���~rąan�Sӧ�Y�e#M7��6\Q����a?A�ۓ/�V=&t�i1X��i?�_2Xq^��c�!�*�4FR.�^.�f&�xux�&����/Ǻ�QS�^v-�6����|�O���}�״�����	���51��y�ė�}�-� h��*f�VȐ�JQ�K�U|q�$�5�*~y1b��z5cW5�]�����k�w�W��9��J�/���2�4���6���0�3�mrYO(<,���@d�JPc�Z�jD�Y�Ǫh{�})�A�|�X#�{�P�%��Z�S�e��/�%.�����r�_��8N�Y��0�ĳ�6e�[:�+6;d��kmo�|�.�QH�0'�1k��Zs������z��x�
K�|�=�ʀI`�͚k掁�S�ÜH�~�r��$�j;��m��g�9�{1_���u�=7�:!�w�`�z9'�Mq؆��fȀ��<��A���%�m8 ���E�+~oJu`�븦�ۿ �s������⺤����ﰌ����o�2���J�<�X@��ݓ&޼>%(�������xb>��KЀ��}!���f�w�ձ���������@��:��/�+M؁r^�U-%��|�z@�8b��*σ��������O�پ�~9	)zAo����*��ë֦�=Ю�^��� ���V���I	B��o��G�\"S�G�����2�;�C�n�4�zR��\0֡�d�d�/D�X�W��[�u���� �(R>?ⷀ��d�u�c�k���4�8<��}w�g�q�
l;�"J�׋��n��|��"���%���}ث��«/�d�15kL{��~K�� _���b.�v��%G8Mʫ\��h\�n��n��L�'V#�T����
�b�"�=��U�By4硣p�C8���Vn�e���י��,G/PR�):��'����"e%$(H���C����mI�
��T��\���Ֆ,3�\�W{3�ft�p�����������*�r�:��/sͤ%�&�2͛�D�'I��ˏTh��C��"���eB˩���`b�H��W��:(��=���艘�NƳE����L�[~�F@c"QC��mt���'ch���L78�!����.�O��+�yX�a���F����]ӰT�p]�x�J}}ݻ�m��̏����Բ����Cmic���{��f|^���vlL(<	��/�'7C��藲�J�!j��n���l��jq4�|��:]���<B��+Fe�V���wh�1_��X��Okp,�������+���IĘ�JVԍ1�K��iE�V�ɌHZ�sNèקkd6����K����\�:�2���ƶ�
d�3!��A1��3³��)_R!�,]
���˶0����f���.��O^DL\����)DW@$���k!�7bt����j��ӏ���2���_r�0x���y�aS�p��	�+ԅO�)e�tnW�yN@�����%�x��5��X�-n8��!���� ��>���w���z���,^`Me�JQy�!��JL�h��2��xE�f&R����%�R�ɦ��?5+\�[�t�
�t�xj�W�g E�W�U�׉*�<�����Z�%Z>v�9�9�a��+��w�Ag�<߉���⩍HX1�0�����������N��4��-1�����B��d�r؆|F�Zqv�2=�a��(�����Q�m������4�c�y�Nj,������SP� oP�I�J:�DHGEc�qL����*��������'U�ޛR#*2YQOȏ<��_�0i���h�S��j�_]]a��	5������P2	r��E��%v-�#Ս��EZ<kcA֘�ٴ敏�w�
Xg$.4j5��?�C��o�&_�1���!A�J��@��L�s���$��������	��J�����L:<C�Ȁ'�$��5��Y���5sD���'���g�RAn��̶M�dƏ/�N>��������\T�/�-y�W�Y[�s�uq��@ms���<"oZւz��u"��h����C:\��Q�=��|�b��ɵ@^�W��J���\�}�{v1/ׇ�̫�l����z���F�d�E\X��ba�\��@�L�>������O\s��05/?u��Һ�R��{Q�D�ry�)�� �[FJ�rbӜ�Ծ���M���b|量I�s���r�v��j}�� Zi���({{G3`���i��5�)�`��Έp>���~u��%�kY�-�}<�~Ԛ7���l(�}(�3�7$����s�?�5�|�ލ��"Zv�VntG�K-f�s��bE�
�4�S��>1O���VS���G&�G�`�?�0~c޳��J���]�G;;3a�ԓ�w×�'����%K�l%�B��g�:�%���!�A���ü���M��*�V���V�ć���^����a�f����U���!���"П��瘚�u5AcF=�e���H߈��u���ӟ�>��o����f�LH��'�4��J7-c����S�H�Ũ��+QP�c�c�)s7k'��~3o �y���\�����m�������5���!)l-��dꑌ�gȉ
��v1f	�"Ղ�Pw7D�i�My��ϷJF�������Q���l���[�Q�&��vɂV$v�l�>o����Smw�by�G��PZ% �u�YvF��3s=�]ĵ�\mر 3B"�cg!�YgI����8�$�x���,:�IwΩ���۝-b�����,�DA�E�tB*�2�E�j\D�(���dm����t�ZF����:w "s�}M���G ���;M���jD[ Oq|�-c����W�r���~u�;�+�D�����T���mSE�[{��'���<d9��]Z�kN �A9�Cҵ(�?��*!� Mo��s~$&� ���yt)ľ���3�mN<�ii}����bY7�;F��ڋ�K/�\UO�*`d`ܡp�	����BQ���<G�P� �V ��"�>�y0���<�*�v�ᮛG�����)�qu�iaT��o~v5cgEu����PŘ�"Mڪ"f���>�;�Rh��Bl��!.���N_�/�u�9�������6�����2��	�VWб�7j�},��\�]�1��D5Ƭfh@	vF`��4��!㰋:��!
8$��~�����A���_�T�����������UY,\X(:����Y2x�΢0�d(Α��U�|��>S��m�H���AW�X��?IM6�E�a�7�[�H�lfo_3$���-�Qr��}%m�ML	e����ƇN~X� E��ebXJu�����`ߎO�l<]D�����+��N��q�e��$Rj{۝���U�����;��(�`!)P8bH��q��s��Շ�6%(���NmmA��o�����o苇r��9V)ݯ��r
��y�P�>(�;;U*�g��I�����S{a�}��#�Z����{3��)�h2܃9�JY��WZ��h�C��z�Z����w��[N�l(;�]�a!�]�&��_6<��k����W��8���%,�eSC=�mV{�xա�2�ҫx� ��vp�&�%��0<��^���ɳ�PʎY���0�x�@*M�MnW �:k��Tj�d0���._[D�dϛ��4���"�e�*���E�'��6=n8�
"�,Wb��.S��p$�B�-�ڽ����|����"ʞ��EmM^���aީҷ~�*ܫ@����sT�B؅�V˴�@+�Ɠ�8�XMzM��$2̨����w��X�56��z|��Z���m�a�<�˲ �����h�q<�	f��"��߶�>�[$I�zg�!����S:�x�{R��$�kp������w!4#u�m�=t���8�akmYK��{���� �Fb�(����z�f#,�W�7����7ygH�:��c���A�9(w,�S���^y�9s����Fh�;A���?����i3�����^i���D�w����.�g��-[����d�1�؃I�ě�)	v1���)��AF'����ˆ���ysD��S��y���b��|���?W8�eh�s���G�C;�T\?��"����M�����Y�S	4��r4�_�L�C���at34يL �i��.Z���}p(���~>��\y�i�7�y�|v>�^(���e~5µ�*/I@ƽz��Nл���/��v̱��������y�B3ݸ���PEv=|�e��
������~P���-�[H�;FJm7�	ZsH,��=g7���σ8%���aQt��;_��2�;7�	d�Z[SӲ�366�k�~$��Z���m�T���/�i�f�� �M�a���)e��%�ł�u��j��j����K�|5UNћ�y�V���B骶��s����i����b@�r܃7 	[
�DYoa\���0X�؁�^�?��+��Xz�%2C9E��0��(�ՄZ���%$ۭ����{��\��#�H�|R��b|���Pf��Y��a-mO��������tZZu\�L�����`Fl����X]�Z�� %�2�^����H!V6�؃��x��b���M��s���gW����"��k�^�\��FK�raY�MūU��9J�
s���8��}�RSkk�ɉ氚�
O��"�Y~�C�]�33��`�����lWx���enyJ�r��`���p]��T��o���Mѣ�����D�}+���; ?n��,����	���h|Xw�xsێ�#��P��U�F�+S�rW�t�X���KF��'�Ip�-�rB �7� �]�n;t�BB#�M~C/V�|�ߓ���6{⤽���(�nr:��$���r(@��F���m�v��.�Iח��`!̫��"ƊfJj�`6,���7�B9���KQқ3��f#��^�(1Lv�M��c�&ǽ���m���MI�I5A�ɑW��W�q�~}n���W=�	�	�G[�j/SC��Z*��W.���W��Jh(��ĸ�.��-!���P��_��3Č���J�'D6$}��lr(m5+��7��
��A��a^�}5���a�ݾ���H���B�#�����ͫ��51�`c�MK/Wt���|ӵ�&,謴��^���7<L��9�)0D= ��'�+�P�����jR��H��-T����{������q�ے{//����R��-�x�c��>�ry��^h��9D=��QuSNKL��5�j�؈IY^�<����s�z33ڛy	�\�m�d�,s�:_�&���'�26WLR4J��GL�$w�F�+�3�v�}��f�Qe�Є:y���u�X"!�{��@�iTѮ�Q[&��9��=M�.ƨ�0 s]�m��Phe�UN�$fiL�<�O�i+����I��OLڧ�K���?�{���C��-c*�)�*ݤ�8\Сy�<���F:�C�y�-y��D� Zv7���t-�%o��G�qNh��K�hh~N �N�4��n��(��:�i��r&�㰨�`�~a���(&�ޘt _RK�1��
?��*�]h�1���]�r�nl�7�|�A�:��D��a�}��~�yU�W&�Rܙ���]c:x�luL���A�m��q�9յs��>3z-�qާn�'􍒾��7&�*^�,�[��ϭRj �]���SL��!:9���}7(
ٖh8E@ᘱ�OG$�Q��skvoB��*;

��{���o�n�U�"6jOVЁ���l�&�v5&����#x0~���|����6��.I�X&H����R\ai���
@�Q2�A�(ǽ��zx�5z,��Y'��O��%���ǖ>�<������;����V��+�P����ϡ폾ix�:����[WǾ���$�>��c|�9��P�r�xe�*��8V��6�6t7!"_����UΕ��L����m�*IYb�aZS#��pI��x�O\��MH/����C����ܢyj5���E�D
�t����9a�B�3��0"A�ލ�/���{�a��+�F2�4U&cV�>�ZZ��"w{��~���Miy��t��[*����ا-���HA?b���&�q͔�~�7c��l��C�o��A���e��i���>��WJ���:ʗV�b����?|����5%�rj�-��k�]q���HKU$����	��,�Z���!�/�.���7��`&� `�=\��<�J�!)(�>}�,�8�U��[1��X����j.���Z"��ܶUA�.�#ص\�Fя��X�a!��$cL�&���~%���%�V#�V��[s�X졷�K��(���kT�����U�Cz��/V�=5S�E��])
�qߨ�Ь��?�������-Gi�jVA�+��?eZUoS ��*�S��e.���GL����x^ߒ��ȟ���	Z��g$��&�:X�o�}3MM2s�?R��Bsw��1݆�<>l��j������ ��{W3��Qj��{�7b�����sS-�H���:���v6�a�s~���^���ŏpQ��mt�)6�NrAFS0�c������B�n���o�fN'��yb,���^<"!�:͢R��F��T�T6�|�K�b���?�q�E�H���^쥇'��~^t�/��x�:�V.�ʱ�˰��/'P��_t���![������e͓f�S�#,~
���fz��s��"�	�Ԥ��.��	#T��-�[�_��y����Z�������a���t7&��%�8��N��|E�]���Of��g�&��i��2�X@�-K�ǩ�����Xa���*��c�Y�$O��ѳ���Er�d��0v<�~v�H���(>����"�7��$�쓦Ƶ}u�8-;+N9�(��=����y��h�zȑ��[�G���f��J�J�})r�誝7��0�9l���� �������}�H�H���k�\{�W�~�����R��d�J���0[��ϙ���51�#x�x����)�S�Rt�ɶ��|�Y�� ~s?���bpW��J6��Q�n��,ga��x!� 1��=訃����::j*�nCv}]�X �j2�'�TZ�����~�M��m�������v�>T�X�j��u��xZ
������Y�����.�� ��!��ɘ�+���帤IKX�T-]�Y��^h(^��YF�7�{'���u\���!��a�¤��K�����$2�'6Td�(��A�r�����I<ߓ4��W�Y�����XQm���| ����#fR�
?����cXo���(��Yg�]��#��7�(���4�"g�rMdKEHx���Ǆ��𡻡3*�b0�u��H�����LH;P�l8�B���5>�M.�y}�q/����hV/H��x�&��8��f�,Y.]�Fd�H� �RC��1���1��}����%��(K����}�}!�V�u�>���轎~
�q��C�
�V{a	G�H��?=R�|JV�-�(B����6�}bZLTA���?�R� ����{�9t�G5-�*��l52�� n)�����d"FG�VK�U:6��bo�ဈ�I�r�{kԆ��O�&�}г�e�ݑH�n���-o i#'����w_��i��(Q)�K�Z��6�����[����G�������*卫�;h~��P[�#=��(��ޓ6|�n�z��������|J���������c#���:X���%����2�6FE�H*�����I��WAz��KYR���R%#�Ge�ъW��w��Iu������ [/�����/����h���/�oB��:"�N��|�`��v��h]_�n��
�Y	4�@JQ�-�Yj��T���C�����ZV��f�%R	A�C���\OB���|TR���W���֟V>���F���S�L�����"��L�D�Z�m��ʺK߼T_�\=�6��C�}L�d���,A��ʠ�wR�B�!vI'�s��m��&%��
~-�Mj����8\�3Q�-�*�:�C���!���s���Y �4�/ ���u�4����Yړ+ǩ���i��Ksvҽ��g`��eE_`���.X+7�����K!���s~����Q2�'�$�>4����p}#b��Qn�8 �9uf�k��J�E���ht���'GTDT`�e�B@?�1���}~Q�	����>I��I\Y�B�̵����綝l�Z�2�����Id(�'�
�
,��ÐP��z��%�<&�,����әz�Q��*�i8�-ٽ�ے�A�$�P�.�T��|�C	��e#Ʈ�K���XǴš�5iC	�4x�Vナkeo�?t�WVT(ư-z���V�r�lŗ��Ғj^��
�ʉ��
�Y8	�2�������*f+Y��H�:�,�r������,��-��*�6�4����a$�u�(��I���Ϗ�s�UEX'�n�� ��3C,6ْjgi�6پ
�fW_8:�s����ىS�D���8/|�����h�:j�$��5H),��>|5}�z�����!�����{��w��OU�G޻m��r�,7-��[
<މb6ԙl�ۛQ�o� ��U\;�=���`��%č&�V��E�P���v��N������1ZC�:ٗ�k�h� 8�~�§{��%�V�u�v".�,󦘑�@G�(���Y�L�!�H)>G�F�:4�c�I�w�K-¼._/����a������G���g��+����
nm�,v�F��m��C�~�-s��;z)a�^��{>Jz�E���W������Y�=�7q+�l)���E�ή9�ϯ�ui��"=�ԑ2���O�R��`���c}�9t�U`�P��_�it ?M`ƜD���U�*Q:W�Fh��F�5�2�/ŜXO��+�h6�����ջ�3�������$����dƦ�B Cpl�y?����<:�g��c.�\h+@ �:�c���������f�6���f�q�@����=�MNQ��Dg����U�\ߛXM�k�'����1u�͠��uGd��N~��Ňg�\�M���LA���!�D���~F:w�er�E���;�g�yHc��͉5c$J�t�]�>ĝ�l*�[��Z��l��� +zAi��z��T��$r��-��3�T��/$��� �b�����/(3Yν��-8�ʿMe6M7�!�C8�7���J���"�c��ZGeS �M��30��D�<Q>�j&b	��8�y��_���w�,���5H�\s�x�w7 M��:q�=���]췭K�V���$�0�<;�C��9�-bx�[�s�������d4#S;��)0B��0�/+���T>�%bG�'�|��J� �w\z��jo�ڏUˠ�ɅG����W@`�H��ė�W1uɒL��a6�`�@ٵ�h��ؗ��j��3�*�4�򥦘�6WZN�0t�G�*zo@Y�٬���ǿU��qL��q[tF7w�A��R#A-)�:g�s96�*f=L��!gK}����7��`[�8�u��
����%�z�F9�����\(������y(���Քc�ݗy���;?�j~6�D�R4h��K-d�:��类޶��D�!T'<� U<l�$l�㳾�"9
�/�����50�LיY,�؟R��$��z�陋�̤Θ��97\�Oc�D�X9��W�L�B��.���u|�l3�tG�#|K�p���R����D��)��\�7�����M��_3���c!r B�t��n�t����p�7()n��'��r���ճ��kY6H�s8��o�]�<�>�fb�uW�ڕ�=��뵣�J��wFQCS�����p�hk];�2� غ o��C]� �-}�ս"�.-f�	�#�2U��ݱ�I��[S���o��f�KGs�������,/�w+��[��K{oU��%�� b�WU[���y���5э�a��=21���tQ|cl�u͠��'�O��d�Wk���9a����t�E\�jI�ϟ��8g�h�˩��2/�j[f�|4Կs��F��GoH�=Ud�s0�-���hG�iH�Do�á���H����~}��>y������#�\O6�Q:�}D�R:\y�4D���/�bj���kj�?���탿nw&͹�f�wo,µ��91a߻ޞL�{����� ؕ�xy��=�oTۡ최%�A��yU�]I
�Id�q,� 4ey�L��Ӯ�Z��>�$�R���,S��t��Ba���[���y$�W-b�O�̥���Q>d꧞D����d�b��`�!�(��=��mm���(�o����b���WF�~6�fT_E|�=Dd���U6������VB�P�k�D�b._�Vbz�}�'2�ի�-�qI�7��>񭤅��u{O��^O�C�b���3ݡQ�-�����E^4���|�`i�NN��g4�.�z��T?���˳v�!ߵS���τ3=��)5}?a���E����ݞ\�� �V�D�l�d�t���*^w���A�v�Y�^L�4� ��>c$�:KD���	�G�y�����3u�"�o��@y����7����:��|�Ӭ�DN9KS��՜�
���=9�r<P���U��ω��{W^�����8�Ζj�OJ�{���a��"MT���8��m��$ʴ�H����{ �Dw7�&�}_N�Z�Xm԰VQ�ʱ��|�ť�)�`��M��SH��@��Sh)J[uˡ�\��v�áܫY�E�G }?O}��n�V�(®la;C���l��Tp�W�Qq�W;0�HI*�c���{�+�I��C��W���@#�H�U���B���F��PЈW�X�Ҫ�?�w	�y��6Ƙx��f�S����6i�BIL�C�{�v�����h�V�27qpKj}�ы�v�	���(C~L� ��WZn<���7#z�1&��U!�F	+�i~�hOB���L�}M�� M���X�z�_�Q�Ns�h-M��� "7Ą��o�p�6T�1n�%��{�H6�mQs�KL�3Q�~������lշZ���5�BxIg��P܆�F��^oC���
ɻL����w�5l����jF�<�X��0���f\�0i�x<C�_��P9(�+��z�`�P�^�'m�&�?l�� n���Pd{E���y�K�p�NT�
��ZTW��2v�>��W����i��Y�/'i��&��?�i�Pp���I���%�ޔ�����|y���N��S.����fw�n��K84/4�����v�����O�Z��Fd#���������d4���Ҹ���Ǖ7`A>��C�L�C/2�	Ɛ��'�?�eB�~���9��I��թɉU;|}��F�J�	�����֟з,4��oWO��o�X���dt�X6�+�IX�B���61lʠ[��� j�("�#����^񘅇_t�6����i��r*�1�\O���p��:�f�-e���tf؉��qZ�m��|ֹj�t�v���-���ԑ>�zp<l���H<ͯ���e,�7T�%k#-|\�f�b��ǜ�j <zj���I��R��a�BM��U���~�֫�Ƴ��@d���������/��0aSn�k����*�~���/T������;���J>C�!A�2<�%1�����ږa�x��b��T�=΁���j�9��x0��F�p���"칑�I�;�S��d��{^%�(�wŶ��ʸdy �L+��$g�yi�?�����R����U��(r� 
3F.[y�q�*�~n������?
����3���h+λ +��:K�FN��4|��Y�;�x1����p0F��ɚ�9����G���d�!�!�wn��p��=��.C��4�a�ZKv���*�`�����Sf�>yLl�ۤ,i����{9u������#�-�#�Z���*SA+� ,@���$n 6i��
���j�`^VE�e屣ᖰv��"kU|��s����Ι��؞�kU�M�g�W`��X�g�A���oW	�|'��-�U�������,�����Q��C��ώx�7O�;ˁ7tT~����k�_�ٯ���!O	iA�
�%�sF棌6�*�rgn��3j�(�0떷D;����O�;J5퀩=J*�Zu^؇CH���,w�+@�I�X�٩i���@y�>�j���8A��NBU26`�~P�,U?������W���|���7}�[��iO�W���D��t87@�~o�eE}#���E�k�o!�J��G�$BP�o[�T��,���w߽Z߽R8�$��,��(�E��9�,�>&�xC#�R談��p" ;�z��|o���bYC����ZA[�ə Ҫ�<��L���߸H�%y-���_*`�W�8A�5���Dn�� ��Q� �yk�,&��6\��5)=���A��<|�_����Ӳ �E�}�<"B�`G~b�<�O�
�wH�{�Բ��Z~� ]�,88`��E�TL���]�<�^HMYEYd���I)��@��/g����l��Qx�+�S��w��>y��-��"��
mũς�����T��˳���d1�UQ�I�J{+U���e�`?��$�ˊ�#��ܑ�.={��iٵ$�C��)�Π;/9lG
�O�ŁMN���1�`�q�Cl�� Z��)�]2H�n?}_9���n��}��_WKm/�����xH�J,8TVIz!�ޭJ��I�u'�O�S��-����%R��PUu&�"<������.l�Xae=do/�F{CoOw	����^J� �"�#v+�\l�vq)�S�;\@��l�uᐰk�teIV�vs
��2���q�0��EJ���-��Ģ$�(�%����8E����S���R�����UO�"�w� ]x�^��QY
kG���冱?��Ҵ��Y�S�}�V�y��W��y5���$|27\b	�So���	r���+aB��C�A[&K�J��I"�J��8�K%�1�Hbr&)_!I�Uc�I��(��%�ƌ{Me�c���'E�sv����w=#�Uܵ����n�A�+Ų{���%T��o5�C1��Ԋ���"�tGA�=�X^1�P+����w�=fX���V� ��<=��TBbՑR��ת6��LZq����qg�Ƈ������<�
K�UX�@mf�$�Z@Y��j1H�C��]�">�����B�h��jQu�˾R��#f˄!��#]>��w�3Ɲ<�V6l�A"�{FH�NxG?+�В�wK��`�ba�b+��zW�ن�G�g��xn�R�{n[�^�p��,��>|7��w��p� �rNi2H��b0�`B/�vԶ��m�!��8-(�]<���[
�l���	�Y��$I%ĘUj!�J/t�#�!I���>��ږ��N����)�w�s�wȊ��w
�헜�\C��!�C����Ր�#��-�"^w��w��M{�9�Y�?t�"�]S�H̎��� ��HĚg��y+|�� J���T�%���w�j� ���|��.��ƽ��y�:D�A�d��햅 ��@�[��lq��-y�@aߝ�WbUgx>R��3�����=��쓱"��M;�xp�2������Y���x�#�zf'���J�2�ex��H�����`��`0��$�� *8�KE;�e��c�ee��HsU�k7}��v�ݩ�B0�Zq4� �/,Ͼ�s<��;g��3ϳ�z�8�m���.���?�	����`;��&�%��]�xnQ^�l!���r�R���Q.�<#��_(;×dhP���&U�K2��<|GL�;m���g�V�gR\�재Foy�����@p��u��E;�,D��Y�Y�c�y�h��ϼ"�O��Ԫ�IM7H�d��6�M"x6Bw��ܕ.
|���J�]�VQƾNѤ�21"���g�]y���[c��@߰
�6�@_~���t��G�%dӽ.e����'�-R�o�:}Hv��}*��g". �T�p��Uw�:l��y�nC�;�:��3:�Ѣw�+�4k%oU�rD�f�8;*Il��ظ�+����p���+�ߛ���
�}�~�U�k�:90
��4���	s�YJ!%[lͺަ�x"�	�Ͳ8xf�;V4�����{����MG���Q͚��>�[�T�����ԃ����hɌQ�J��L���#0p�����*˪�/x��$��ϙqnP��մU7  8�IDAT :���x"��ì�Q~�� ��M��{b�Yv��}��N�5���[�����n&�M�du .�lxM��R�jE8���ݒ���~̘~ɵs��=��mK�4?;�
ޭ�v@��$84� �;2�n�tc��Y�Ņ��¶�5po)0Q���,$���w�w�̈́�
g�T6�[+�0e��qm���sl�q�[T���xE�Z<�)�h��Q���1|!�	T�͏LG�������zĔ:H�;l�Q�{�f�]���<w����G�R/�?���j�u�=Op���v����l+���� ������j�H�R�,y'�5�����~Vf��d����H��w>��T�`�}'�ŦA=4j:��i��W��Q�Z0�AuLg"���
�1�j}��վ��2�4�m�O�|�	�F��'".|��Q����լ`�}8����&oim�te���G��
��c�F�|�J�#�UR�?��t%�@�p����.andIi�:���}}�V���g��Ԛ"~-5Hnl|�,n8J�P��S��X�DO��B����J<����p��wj�Z�>���X�	�m4|o6dr�QX�Y҆-k;��s�0�-o��p$��	�k��z�8<5P���l:�^3$L�o�SI�:�!�)%��b��yՋ��
�b�,Ր<%�5�TY�=x�3t��D��dс�{�=�
���i6�e��+����PJ�eo��y5�YyL<��(E���o'C��w-5H���%7�x��/����Z�YbI�� �P�΢y����9���
�%x� �FO�7� �S�w"- ��z3���F��<l<"��J+�[�d���B�롍g�f�_=�P�#͌*�Uom���Ha��YӸV��i p4VY���U�g�[a���d�������']�/�ڨ'с�<ū��7HR��r�Y��ƵFlR��W�Ӽ�+
c���*p�yIKJ9D�eyP>�1������/A���L�;���$S���$��!��P�/��e��ߨ�0����9<�{]��c��2>,�Urt��^ob�륳��@���$-!�*�R��~ xg��r3���9� j��� R ���'�J)$��k�z-�y/_Q�z�.PI�q'��]���
����e�2�^�0�Z��b߭l������©�i%4�A���t�p
�YyiIһ�i�;;�g�l�����n�	��cg>z�Rd�m��+l�46;
x�56�EZ0sA܌�����p/k�=�T�O�����L�^A$`�:��w+��w����hۥ���.H�BR���E)W��q��!�ӎ��o���@�)�*]o4JƸ���x�七�Ѭw�1H�1��5y�
g���N7u�g}�P�w@��C}]aP^��+��4�����0����N0]7Pi����Qc�+��})FY?f	�d�'���~[�181�(9��g��D�֢�Ģ���4d���D�U���15Ϊ�#�q�류�,��Ȍ^��b�hŴ#��wL�T�y\�}�4H1��C?X�Y�w�<+���+b�1����|�ʵ��3v~J
��l�m�����w�ƾ�3�M���<��`��%$�M�-F���^x��c�+3F�"���`0��zv�L}N��ژr��5�3�^6�(�+D �,�ɫM����נk��m3�}�)/ڡ�)��1LT�����!�C��fL���
�^!���T�����y�D�K�t���z�$ke�ݑ:��ot
�B$�a��5�?�$�{�� �Ĭ�h"ć�*�ag�&E4�����<���
>|W��\~�W���`ӭ[		��,1�u�n'c�1�`�Z�z��O�!�3Buӑ�NP݃)z}0=��5��4?�5zd�,%/��ƚ&�ۚd=X�=��qO����28P�J$#]Z[�i��1�7��a+�E�����SaZ{J�f�?YW;��wxK�K^ذ*Ɲ�m4H3��7��J�4Hy��
���I���5�Dw�|*?�[@g���pz�������g3��Տ}w�B�M�+6݆�t߽��W��Z����cÍR%�β{��H��ČU]��k~�t;��FRhD16�fA4���J�C�?<A$�;c�I�z|�}��f&'�;����$ߝ����4���`ޙǫU�ܑ�(��͡~������<|�=�&"��a�8AxL��1�7���ee��Щ0M�ȳ[��*�5I)�1��'�����N����p鱪��R�fµG���MG	�e/!�je��ӽT�1"(��FNp�c�O��M'����ױ�tM�^q�p���ס�ݾ6���AB��{�_q7�RTT�jjP�����df��
�Z��m��1��Jx��U� =H�#�{Q^t��uY�~Pp��R���%ם��P�N�|�}O�_�/8^�\F���7��l�2b���]#^��#ke�%1�QJ6�(�A�p�໬�,5��+p����`�@x(����@E�x���U����*+@�2 >�s��&���B@v$��]'���t�����W��_��[0���Ö�:�m+a::��� n/�r¦�I7N��s��չ���(�����>C�r���S2L�J�c��+5�m��5�\y�����Jt�dt���[fH��*�3_h*ߝ��W�;J��=�4�o��[d�!_�!�~m���K����N�=�E�(�����O���ȣ�)�T(�J�'�gW���j�R�E@�+��;=ߑ*�ݐ6��VF�oO��5�;]�`��t�-�A��$�G$��Ȁ^��0ݞ���G���t߿]��Wd7�^�~mC���S#��/Ť���FŦ,��|\f+Ն�M�/���i2��nKF����M�9huL����7S�3^�yMI0Z�*/��+�SbOiA{+$%}'Y���F7N>�?�?�I�=1�6��V<�1H��ze1�ë9��l/�j��퐍<�� ���d�+4�*���
��L#5w�wgI��WU��=X�d�w������gY�����+��(�Az�^R���W��)��ږ���V���׌yo��.��X}�>7/�=���	O���$�E��򗶤t:@Wl�o�\æ�n�l��Rڨ�둇$�|��T">ڃY�n���	�#>�x�;Rޫ����d���Z�k`��*��'au�6^�0u�ߺ��V�]�e��0�V%��	Fy�o�7�O�ѿe�$�#�s���Z[$:?N�ξ;0��J?�u�c�Ln\9<�0����*>�#+O�w:����-|��٫��>�E���C��A�|Ħ`�͝#cS�ؠ,���GZr�K��'�$b��?��G
v}$H���E+!�Ŵ:q<�N���:V�,�Dۭf�e�őq".�bs$��`�;���$�t@zh��M��sF	IuYc�I��_�XAEY�
7��5���.�(3����$�����m�� �=��H`���OKj�V�C�|���죭����L���L�C�}��O��l��Oc���Cu�$�]�G�L��/A�+�P,�W�Z�Q��s~,�a�gTyU{&�讒�ޝT�WI�5_i^�'��p~y�2 ;�8�+�'��O^�6ft���VĎLؓ����t�5�1HT�E-\��Ȫ���,���Dn�aL����3B�)�x��J��(YD��h��$���]$yH���� E�\�JW�}��<�UR��w�Zk�٤�����Y�����C�*�>U�
&�g��
��V�ՓBiv1�n���^/+��JЫ=��Ķa��ֳ�|�f"2����Ց�Pqf��V�W�h�l<� ��Q�i�P�_B}��T`���3��.ZzYH2&�J^�iO	�����z����Pd��C��y���l��<a�!������$#�,	I%c6pz�25�
�C���	Q��JRЯV�,s�s���icN��x�\+��G�$�Ľ���=��u5�4K���r�9C�7���z���3�Ov�<x��*�*���&Ɂ�D��)[A�;[���+�gtuю��h��M�K��l�mAxƦ������pą�uN��aP�
k�F�J�ӊp��gb��|y���cL���I�&\�8�LV�z�H�E�.3N�ƾ�3�

4�l�n-� @��O��r\�n+��J�ud�k�u��BS1?2h��ƕ���+eD	D�b�6���~ϟ�gFIrr�K�#!��A��h[���a����~V�,����4��̈�̤����Y`�?(�]��]�$�tkZ�QBB.l:�_��b+��#.x>E��?�B���ݎZ	r�^g����(���@�y�Q��Qj�j���+�&i&l��R𬌏E��({�Q�E/��~����=ɪg��[$h���H�+uN-l4����Pq��l�E�
=��9���_E������0Ü��I�b�Ӓ2	Y��
��f��}|�ImM�݊�X�=Q���z����%���ʳ_އ*�&i%	<s�]� ��A26���p6�K�r0�^�|�In:����=�n����Ԉ����>SQFJ������A��"�:��Ѷ�Ǎ�n�e0�	k�t����}��w;��o��%\+����0 V^�u��E;�O5Q#�K2Ɲ�G��I���P5|gz�N�wD�����VI��k�I�d|K�	邅���V�u��R$YI
]�W�>:� �L�Qu�
���QW	��ɁY��'N���g���)0(�k#���*�>�	�T���J�ġ7�8�h�"L�!6������Qg0��zՅ��;=6X���t�t�,	<���t
z헧�LW�J���1v�� `� 8�cT	��F�	���� ��-MX����^M\��톳,���~�Z�3"�z�0=I��nm�\��/w1�m�<4C�sy�dn`mDDd���5��������`,�K�h��6��Ņ`�ƶ�A�`���0HQ),�1�N��/+�?�=_����+�Fk��[g���<�nt@�������7�L�o�L�o���,��B��º��!�%o��W���t�#�.i]����N�J����|�3�y�+�z���D�� 8�uH�H��4U�������.g���g�ZAb�Q{��ZM��"1`I��E<&yKU1�2}b� z���8R8�]��VԎ�)VW�����-������v�~ݻ�����wǢ}	�}KW(��I�wxpVy����}G{
|�����[�"[Ij m��[�A:�_(XЫrӽX����t���tŀ�� �t+��=>2s��|�Uz���YD�.�n�y�w�l�8e��W���}?�/�D1��|��,����D���d^�on�_c�,����Ҹ6�/�F��"��a��4`�*�@���FuY�w��G��+V�cY�ob��������I�I�<��&%��}$C�x�~C2St�A:����g߽�N�^4\v�������9���yŰ�g�����Ҥ���*����s	~����rٝ�"�ukOM0ݏ�d#2�tEd��T'c��W�C`:�C9�0P}��(mli��,C��`���
|�/��S,*�����d�8I�^1��=c��'i��c|�`g����@�5�.|�۶��T{*�Z�����D|����N��=\{�_{��F&�"P�-o�⑐+k��+�ĸ �F����MZL��⒌M��*�}���;� ŋ���U�1�އ��}�l�IE�<��Ϛ }|�@6�|'��O���wE1HG:ot�A�v:��rF�G���Z���I�t����h=LGΉ����/x�W��攉a�h�*!����$u�-�{�b�)��$S�&2��[jd(8,�%`��Ar�t��	�	L��h\F�$��RỼQ�m����<�ì�,�p�HGe�u�H���,\�o���,ʹ3"�A`��$c�P%IJ�cliV�0#;�QIM/w�AB�����;�gW�U��S�EMj�ߛ�u's�Ĳd��h�k��{c<��f+`�<7+=��ľ�D��Ӏ�P)��`ow �{EЫ�t/��f�%$��y�G�z�O�^{�Fn�ϕ{In��A6�����2�� �bB�=yJ1mС��#M�G���|��'��}�l\��+ig�����~KN`�loi�ļ+b�1I�[\Q���Q�o�*OO1��w>qs���Nĭ:�aG���|+�TM��
�iA�
��l�zy�m��d��I�,�ga�<k�g��� �l`�"��ȟ��R���b3c}j&��bL�Yhuy� O$��qVau�Uo�6e@��TgI�Ïnp��~�|Z���v�����n���N17�����t,��0�E��؈��{[��+�3R+N�9����w�30���3����^��|b��|KOi"�|����݆eC�F�����肶�"8�o5V4dk ^iy����l���X}�*K�891���1�$9�P1H0		��Y���
����4I~���f���7K��К;�OT����/�;��� �����Av�ʳ���h�Gy�Ļg�N$��e]��F�S�\lF���X��ƝY^;=/i���#-N0�\���|l��Q-�ʢ�0�x�}m_�IǍS�&<�8Q�����xU���_�S��Z�g��o19#l/)�)e�R#������Ƶ˃�l�ɡ=�%#ҍof� W����R�\����厓1;l�+�+m��0l���`�/�<��/W5A�mb����)���C���҉�Ϛ���d�6T��*�~�p"��!�a�_5�D���~1��EyJ�f�&Փ���M�1>��>��xlm��8�����
��ui�00��V
�zF��^�
�����������:� �3�I��M��Ԑ@z�J6����-*<K6��c���J%}��;��@
M��S��:�6��H�P��=��#�0-�Â�|q{�md��9<\���VqU��U��m2:�|��Ӓ�\��A���Gř�I������qs���ij�e�j~��U����Y$&p��"�wv�6kj��m�+�R����Ny0�d�0H4���c�T��Tg��^�o^m�|t��
t=��W�y��@�����t�V= ��5��s򂌴 �(c�QJ��MW�o.�{��bF�Kz[\����
ڱ.o8Oj���#	��JF���w�%ȇ�� V�� 5��Y��_)�E�WCW��^4���
�Sаe7	 ٪�s�� �!�-I��T�O�Q�֧vW�v�O:��\�o�A�+h��Y��9����W����� ZˉW�ʳ~��׬^��F���[Ҿ�W�!�Dk�A�����0F�X����>ц��6�8�I?c�2�����e�$���x���P���ȦSF��@v�'��
�Dj!R�j�oec�'4t'V�:+�J��F���I��<����U�#�wxJ�Q�1\՜g�R*ue{�VO(c�U��F��Jo����Ƕ->TzC�!�,w�?���+[Cdݕ{-��H�dL6M>�t~x�~ȕ�XV���f��w��n��*����~�`0�(_����Z�~�?_�j�+�k�l��nP�Ā�u;���%��Kb���̓��[��)��`:�^�36]Ӎ��B��t.���}/[@ih�$h=P��=�;�M��:_��*�4���#���7�-<ۇ`��'D&���/�
��vx�����.,5�p�.��yr���U*��^#`��^�Tk�H,܇�o��2H6oj�ݗQ"�P=��F$[	�>B.��F����`ϕ��9�;��&-MXE��I[�
���+� �y�w�W��@T�W*��Ar��Ь�[����5���dq`�--���ܬ��'�`W+"����G�������l�3W�Bt`O�\Gc_iM��uI��Q����I����%�h�Z��M�Y��h���$d�e�M�L�Ug7��^��o��*z�&�V��kA�6�n,+�#��GEc��G��H��'a߂��K<��� ZZ�w����c`0����$2�w[R�%&�L��U���F)���ܘ�ܣ���7;�?��xЫXf��nD��bn�A�{�QBB�B�n+W��R�y3x4j%�$��S��`�-cQ�7=ݺ���D	Wy؊Zc�յOlsFp��&�"%�A��L�+�Vy�V��H��B���
���d���캪��s�q�a�ŵ��1]��n�A�!�Q��;1�ǳN�,�b�1��L�񓭐>�ƽ�̀J!Pa@pӾҿ�7&���b�⪴Y)n�I��)��:E��H`O��"a�=�'�UA���P����K�G��<&0ya�/�L��y厧�ȹ)����T��$����[pc\�ĝ�n�/� !�rdBo�q��ؐ����^�C��8q=�����93H�0�7� ���Ho#������(_|�{��Ѫt�w��9�����kE�-bh��yK|���I��� �ŇNIu^*�WDN�ӕ��B9�<㎒(J{�7��f�HW�}s� ��Tb�4LŠK�"�L�.I%��(�vm��
<$�F1�X�����W�S��^�`�K�����<?���{��7O�\���yw�7� љ6���PF�_f�g�X�ʳL�R>0^��V�H7@���e1Χ���|&���W<�H�A�7���KL@L�F���u��9<β?(��Vؗ�wy�d���d�@Zq_���4�oy
8�V����p��6�R�Jq�C��ثI\b�Zu���W��,	�I�1H��"���d�����(�����Aʍ�9���?�X��U���-��!�[���G� �$=��>��FZ^:u���I�4�$7]1KH��(��
-�a������Cn����/��Abu[��6ʵ�Y[@A�G��p��~&]�$��JÓ L�e��/
�Nы@)�tȂ�-�tN8��:��嵲^�Q2�O�x~|��QDJ!E�} �����Aʍ���|��ٷb�!U�,%�i+R�l���38��<7��t�R���t��Ķ�rӝ�����0�J�XquU�]���W�����Mpv��g���[6�ݝQ!Mp챴z��'��F�TB�퀼��h�宑�0�`���Ғ抭U����_���*��d=��>��g�!2��d���d����^ٳ�7����~Y���7�� ֑���XM�-�Ie�����S�W�<�DZ �5�t䦛�r�%�����A����:l�{�AxU�w6�1	
ښ��jc�D�Y�*��`_�#T<^a)�T�R�R�{��3x|�H��od���WR֢�,w��Ir
~�T�U&�Lϯz$�TFs��V� a�Qj��Zd��JW�OU���M� 7���V��36����
vu�n��tV���֫C��Ŧ��Q�U�[�v~�.��@�Opl��@r��o�5�V�N�
�s*&�x,�I�4�όRf����|4�:I��U+鞿���\����"!6�y2d�!�"�"����b�����Ft?Ž1��^co,�2]j��&5䂂g-���/b����Y��'i�C���@�'S�P|11��?��H�������}$^ob�k�z*�x��f ��*��j���s�]�$�6�����[�}ڬ�Ʉ~�Ϲ�h��|��e�eWUqU�"@<AΞJ�����ĲV!���@�� ��Xv_���e�_�a��7[<�����w�D�� ����3n��=�����J��h���ʳʁ��ivz?����:���Ց�]���g*Q
z%7]��4I�bee���i������o��C-������E?��bZ�s�����}��Y�Y7��.��Z�A2�M���
�}(I�>L�V���Jo���H�)y�y���ͮE}��Q�
0�� I���u�� �5]�y�����YS ��`ߑ<�N�x+yKi�+�̺�������T".��nʎS��t	��{��~����,�o5a����R�[�g�������H q�n��Mm(/�����j�d�����Aڀ��l�K��fIu��+�J�l����W��\�=Z���~�͓A�k��s���4�l�@�
IJV8O�+�D@jbߕQb�_�E��N�:��G��cU�}<3IZI��5�'�M"��}%&�%m�/(M)���*EO��w�XU蘍��������z�G+dH�wݗoD�~��y�<T���A����ԑ*}�+�O��H��6��Mڞ�Ep�-���,�b{CV���� Uٛ��Y��#5ρ`!JV�-����Qb�U�����+����ugtWA��!)�,���4q$����g�́���^}v}cS�X7���ĝ����ܑ���q���Im�[f�3�J��2�/�J#Hv�e^��E��$��P�I�sZ+����oR�7��T�U��ջ�F2H��2�;4$�T��J=|G�YI
ϭ
���gͭջN;�e�4�\��?}a=!����]b���W}�qAu�í�Dj��6� pϖ�Y��}��^D%Oˍ�� ㎴BH
�YkaJ�<����AF��M
�չ�3N���4�6�c�Ԯ�L��p��A�`��^YYyK�S���[����b·G�6��5�xr� ը0&B��$x���L������{��1?��[>�*1!L�s�NA�bё�����t��4pKH\���!���>���X@dK���\����wڣ�Lw��.��:|���Ӆ�NJ��*�3q&O��>+/	y��&�~�:�7"�rq�c��	r���a�l�� =~pߤ3�+��KK�jU�~#}��t�b���ϯk�-�v�`=�^)x��ή�/�?Zu*�ط,�ڱnp�/>W����h�tw�q4!�N7D��Ħ���k�t�$�Ķ�M�b��Ja'�>^��Բw���u���m��6`h�԰`��}c������N���rf�@T:�z0Ӯ�
��I���Z@Tc�X@|T�>�O?y� `��WeE&�t��<;���)�vC%+([�� ���k�k��M��$�{~gԑ���מ�t��2H�s	�+�xy����-���1��;�[>q��|���Y�UJ�io��Uڋ�y@��.M%Y�һUQ�9���4Xis�`�]�:ͣ�?�TH�E� �9Yͫ1H,2̫���F��_Uk��d��ћξ�
A�[�gW	��/���.�w�P�A�د�`׬���Wz%?�<�|z���i�/�wd�;1�|_I{K;��'q��n�U:U3Z�W,G&p�&��Zu��ƶ��&��W�C��u�L�@�ο̴����a,�K {������v2L1�YˑR-ں�B�t|l�� <�h���U�wk�+��.�w(��|��WQ�U����<7ݨ^a�yn:+��.�t5k���g7��+�l��Ƹ#@��8:�;�*�ު�TJ��5cJ*�PY��;Q��o���=��"�2��!M��+��_�(U[)�!9�A�]O��¡�#�Z�Uὧ�;��8K�u��s ^?0�O���je�T����C�Ҟ�����jw�����/JA���kB,致�u-�6�{Gg�Z�א�� 3 k�J���:NZѤI#�Re������H$�A���_�Q�K���Ğ�S5��|Q����ɲO�ȜR�:�|G�Փ�Y��@��zV~'6?�����5�͔�^e��M��F���Wz��^��h�tBV�A+��N���a�;�8�A���==I�	���T�ު��}�ڑФ=��jU�x���a���lϥ�{cdk?VP��[�Vm~ʌd9=�>BޟS��̋��F/9	�j9�A�E[�k����`��`�����G�����!��1q�^d:�0Mf/�rz�z�\^#�aV���t��L��aq�3�1�T�F�5e7pf�%�;1Xl��B��"UibvZ�c	�����[RV��E���ٺ�������	��j��l 	���(�9V:��A"u��Y'h�Q�*���A���+�-�wl���Ś�Ϊ�����{6��z$S�T���*�{s�#z�z2�����t��n|(�tg�W�3az �g�UU�@��i�T\T%RU]��&��
�]'��u��K^;5v^��㭪2H6�}�G��4����f�5�}�A��}��䕎�A�S:$`U��~��"�Z�d�j�V����A�}��ވ��jy;�\�	/�w�b$��3�,�F������{�@�RQ����~�MGЫ�t���.��
=��-â����P�E�j|��%��t�Rl2�&oK@�CY
U\e%.h٪#B��  �ӮZ�t^'� �!�}�6�ȟO􎐼�\f�P��)�3�	c�a��H�mU�^[Sd7�.Н���
��;�/V��]�]Z�ZYuzU��������p�&]b�]���9Nh�e�މ�ܥ����̴�>�k��-&q6�[$���HK#�}d5{b,��4v�U}$��:x��#�Q� �=�rC�A��:M�X�a�G�AB�r$�T�����<|�/���5�}���wk�*]!���,���������{U�&��P�g妣��3�!ǆ{��`�dm����9s�I��� ���O˨����Z�iQ�ɸa��yR����+1��}�u_�D �M�|������Cg�+:�l��.�Ԫ�Ab_��-w�e�|���N�>*���;B�r$�T����^��q}�{+��R�݋E�w
��ME�;�3����0LRJ�J�xgy ���2��0�.�M7���)��
� �*�F"O��,�o��lF��2/@3�t�_o�!�D�
�tCuA�m�/���J��E��U��W���j���tO�{2L�+�����c����oҘ��Z0�WM��k9�A�E[Wx/S.��x?	��+�4���SA���������=�7�A��3��NiI.��򿔞Cd3���\�^�*�x� �����K��y�0 1���Wi���c�������WUAvy���̴�#}$ ��"[u�j�b� �grLH�	1!���)�!YˑR-ں�{/��{�!�� �e�g���߹A2�ή9h�����g��-���VBb0�����k��a��Qq52�,Ai�I<c=!����US�\W���a�h����i
��pf�u�%��|Y�U���Y�I��$�NCb�&�UJ#3HQ��V#�A�FKuzO����۳ʳ@w��,��L�A��<�TyUbTXu����9��:��tu�����L#U�댕<&K���'>2<���@D ��M&�<6��0D?g��횽+�k�=$g�M[u\iWa�ճGa�$^Le�hG�A��	�}#	�/)�zvI�+��)�������l�s����TЫ�9u���S���	�^�#�W��76��ͥ5�L#��I������y��  �`��)�Y�}`�8�A2�ʹ�M�)�Tf�k}cI�72J���n���� :
NČ���Z�,yH�h���e,�_����]	Y�.�t�N���;�� �����!Qj�Mg�#R�W��g�� ���Iz���d�EV�4�AL��@��=��I�+�$�V0Dϳ}$.#*�_t��4}�T� 4�V�D�ƈ��=+I!�U���ӝ�ɯy|d��w+��(�r$�T����^�VL��W������zuۂga߽$xV7�� �@V��;��=��*�N
 ���{��ב�n@e$�j�l
M��@��F�7Ho}���S��O��� @+�F���ו�R�Z���B~�IIije����U^��A��<4ov�v"��d��p�A�J���3����?
ގ�K�S�c:��ڑ��s2:�Y���L�5�*�7J�Zn:��TPϚ��J�^3��<�Ħkd�4����4Rl(�$�r'���g�235�� L�]Ԑ�:`�a���g$;�;���G���Qw���7A��Z��r�s�ׯc����j�x~3J!���H�m5�l���7DɊ(��?D�	t��wѺ7��݂g� q�<C�a�g����z�	�k�(k���'k3F�yis3V��y�T� �r�s��-!��騆���}W~?�=#KmZF�Uǵ��2��N�l�Z�&�Ԫ���n�}�fUy�Vv��n�����ỌM'kDʔ��
������y�WAu�bԥ��4��g����ZҴ�[&38����.��"�X�'U��az�}�}?�}���d�eוR9եכ��!48�;��a��!<2��/��; �+��t#~n0]d��MGЫ��L׌׺߈{+�[ѳ�� �a�����Z0��JA�0źBP��'�9�i�e�t�}�r�s��[�!�_   ���j��  @ IDAT�yc�������Z��d�$�����罹�9'���$��-o��]��>�B��d�"%�ݤ��(�lv�Q�OU����R+�>~���?}r?~v�|��������f����m����wﳻ�3��?n�X�]��߃��]��{&�8�~�8�~�0�Ƈ{��P�d_��$�Z�5���{���{-������d��Y�ŧϟrbt�M����:2�����vyٽ���}��N�����y��a��ݹ��!724$9�&����ĄɊn�>���++����;:95yO��2n�:�Ã�nh��I>��t��L����=(���¿�p|��Ϲ[��ƑɟV��O��+�f�������>ڵ8�����3�tf�=�����n�.7��]�Q��:Ao4y/e��&��W���3H��vc2D#2JE1H�kkn�$yxt�e����%�T�������@8���V(������׏��?~\�\�!*�)�t���~&o����s�n~rPr�u=�/����ti�4�W�.��1£��U��!Rt-�#�ntH]�����[� I��cu��!]���⏧����'���Wݟ������+mg��?~r_͍����e�0FS�!oZ��� ��kN��B$yG���Cw �h_2�;���K�98q;����ݫMg��f6��d�� ���77�.�B���<j��9r����K�t�A����ٱ'V<��<�d�:��U-kie�P{H��������{Z�����[Oj��q���nX{E�<�p�y:�y2�<\'��]jwG��������A�;�`MWz&x�\rim߽Y�sK�{��֑{/��^$�\�.S{8�3����uw�W�~�x��/%�d�El��J�]MwHg�	v]�Ʋ�Y��A��59�n\rL{/#n\��Yv�=$]�T�,����l�]�C�t?ޙ��
��=<q�g�O˻��nO?�����K���)<��AF`x45���D����ݙۼd�J��k�*��	�l↥CÔW��ۈ��Df�k��c`�$�j�e�����+��tG��GѼ_��M�TpO	oCTV�yu�92��F��I��ј���	�%�%����������2F�S��M�@�V�2�V�A�Xv������'0H���y���������`�!����L�f��-�X���e�-�h�.*�[�R��;�72F�<0؎x����Wz���O!��!")$W��=�#�.�|9�����y�70C`lM�~� M�*@\0�8A�2Fȼ���a::>qǧ'&�.���{K0ݡ`:�W�t��n[�egP��r-��o2�Sl�Wrss-���C���a���/�NÛJF�����`��CP,c��
몓�z��1#c43� �`H	�W�A��Ou]�ol\���^��~L)���@�[����(�K��v�J�Ctd:`b�UJ�����b�a]��^���R)}^ӯ�1q�P�1J�u���?fv�]�$N�f����h�� �>�69(c4���y��D������ ��TAxzS�c/��WK)/����1��M��`�ѭ��D'x�I���O�K_����%��~�DTp(ᢃ�{��w��w�H�w-ggdcP�7�z#��%$��f���u����vs�YyI2F�}}&�;�ƽ���۷e�1�#���A�9�&�(��O�W��A|�.��5XU���r�գ����טM�Ząׂ���OL�!��i1:%I�Q�<��}`�ݣ�A�H0����@��x��}���SwrJ�Q$"KH*�@��#��8;��gg���q����O=��1������yzY�]���T��c��$���nBaO��]���â[&�u�P�����36�\~MԸ�����6�4�rx�����@���uj2�v��*xV�������4�໦EKz|r�N�=�D��ٱ��+����ZxU���䪏��ܣ�y�X����z�d^��˥%3J�z�Y�l[m-P�;�C��.Bqa3�����R�bc����Z������ެ�(���9�te��ʝ��so�W���ϟ�Y"Y�bf�IH��o�M��=�rߪ�w?0hx���n�	�#6Yd�>&{�:,�P������{Z�HVjL����/,�'Yǳ~��ev��6�����/��A�(qf`�x{��4���錠Q� �w���b�ı<Z��&���ӏ�_`N`��M@e�1�^o�r2H�v���nOA�;���Wl��9�V�2L��T~@�|�-:<���� n���۟͌�gs*Q�pԑov���*sV�}ע�i������Cy�Սu�����6�_k�p��Oܳ�E�E����o���[�p����� ;3H:��Ռ��d�A���7c�(�x�b?����N�w��c{Q-��3S�#�hd�(ȋ���S2H���пL�@�9�|Ы���5!mR��4�=����YgB��ԑ��B��E�:m_��C��S���u;{�'U���r��n}k�&����c���#�T���:����bTl/T��{Hoޖ���R�ČY4fD��A�@��b:�թ�Q�Yi>���	��yH�3J)�Q���s�+P��t"0 ���+�t�Ǧ���+�ľ��0�1��$����}�w���6'���+u�����v����-�����5@v�� �b�ԑy��ލAz%c�Cd�S�A��1�IcN4�<����=6������<D*�"m/I��QyK���!գ����¨;�A�2F�ۆI'�nK0A��Ȧ�W]~���.��?4��8���I����S+�Vϑ�sM}�Nuv��ą�����wfoQL�l���<��/���?� X�2X�[?��b�b�bAl�řY7?�c�`7�C}��A�~��U���ӓn�=1Q���[�3�*�������I�+�f��>���GI�CV�����F[�%=j�wcC=nLy�F<���Q��G�	�k��x�l��A�s1�Dp�D���z�w�Ŧ[�{Q�Wc_�x*������5$&z� \���b>�̋1{B�W��d��dE5����~�CA�dѰ�0A��f�H���o�36�ᐯ��^ݵK�M��o5�,�
���g�Ο�+�}��Mي��G�������JWP�����w�ͨpz��J9��Ć9�H�g�������$�H�W�k K`,�.��y5���0L�d��,+���r����ׅ��ļ�9�́1��)�.�#���׬�c��h��e���,'�Ԅ;z6��̼��Vv%�	����t�Uaf����p+�'*8�+�����g%�:��*����C���� ���~x��F
�}M�~��!�Ж�$B�%��B�˫�ABBa��{��Z�A
=���?އ�.�!��k����w$�}+�ߟ��|�F'$��	X�${���zZ2H�h����*�uEU^����A�tDǦ}��h���~���Mm�!�Ruvh�ˊ�}�x�r�%�]�X��e���^�[<	yGtkٖ����[i��w5e��2B�HB��]�Y��*
�&� �]����3���O�a�{���H�Ð��%�B6)�������b� ��ӒA�G[U�kL���Xn��=����
v��]zMl�*jԟ.$��wr���+빠Ng�|Rrҳ����3v�ǱRk�,�R�DH�3�I�]^)M�ռ�x�k��D#������ە\��R�pk��L�\3��yD�eA��<�z�$<$����Z��^�+��nA��z3h$�T��Uy/,:`�]���r��[^�1��O��tUx�O�R<k�K�ZI>Uيg�CD�g��|wA������+/"L�kbڭ)���ĭ�Hg']��l���h���瘿nK��M����E]���^� �Q`�5R���pzvj�a�B����� ��e`1H�"���d���V����[LG�M��20 ���U|����<�T�@�O5�'*\����uG銱����.¾�(��B��*0���  v� Xu�
�{������[̬+�d���8�k�"�&��{n��k¸�뒧�yK�0��ȿ'B�bf�	�ʫ�d�G���Io�5Hą=}�3h�}_���i� գ�K�=���6r)�M���&6�%����l�律�w$b���w�Q��~=�}���.�w�P�?�!�!�I��*�f�U!���K��M0BH[z؞��-�v���B�,�AI�1��o����~�⪪_�gֱ�bY�{<��z�v��@�G�5�~�<v>�]=���O�9����Q2H��[L��^��V�5x�Q�"݂^/�o�w���HR��:�������*�R}v�r��N(��r�yh���aŵ���*1�u���I����B���)�!]<�� /6��0g����_<TS�:�u+6������+�="#��D�Ym�Y���cP��%Y8+�A����C�Y�3d�{�t�1J��-0l�eI��*6�	��u�Mw�V�(kpz؇���A�
����h�磌����H+3!�7��9;���b���'�p�jI�;���d������5�gcj��`Xr��5�z+^���MF�z�*hT�j���[2�Sp_�]�1(�V�4j1H~q�=�����%�T�] m;�.��NL�%��TyU���ꁕP �JXjMӀ�o=�U�4�N���
�����;��Y���5m.8@@�@�1xWT^q;��R�Q�-*�^>���̹ѐ�F{����V+�z�S���Y��ى�")i^-&�@8Y_�p���$xC�R��[�L�λ �n�س�^A�G����y��ĦNz��Oo�C6=dF�R�"�g�#���d���;���ա�����[d�V'����Ȋ̺�[� e�VH�IҨM�#&����eH��
Y��S���tB��D�:ߋSe�nE8AZ�[e`�:^��r��B�A#�@>Q�iK�N��0%$^�ޑgӝAp�M�c�j`�Z�5�a*�:��FUqv��w��Tي_.NX�
�HH�f���AAl���lE]�$b�����Rپ{/�y��i��:a��5�z0HH ��QQ>����B�--XH�L�1!-�`79�܂��n�c0��ˮ�	F���)7�L:~N0]Jl�[�*��w�#��TCT��t�UG�+p���	�k�h0�Z�@�_L�^��N�_Q��j9�.�I�X ��r峹%�'��5z���Уmo,�"=bU�Ж��h���(9�m]��ء����[vh�aQ}ya^,^�Ɗ�@��S��y��4�C�-�A�Ae��N0��ѹ :1��SЫ�M�K0]Jl�[l�!�z�gs��L�dfX����\�<K�̃E�v{��F�bh-k�[�^��Oʑf���9�0>@^4�T�@D�,7��$�,<t������#��鿲�딴��:�O�w�#}���(�dp�;7���?e�ؐ\L�}1�`��b���M�[I�iPhpF�-�4�a�#��s�^~�A�@u���z2b��j��ç�4H~J���d,Fż�}7*�/���U�M�]���&T�%�us[Y��L�1�������Vܘ%K�	�N�n���P�mA�Q��/�mfY'�y�GV��+YJ�#�+d3@��Jvy�V$�d^�A�p�'$�}(c��iK���J0�6X}Ы/!�.�M��t�F��Aӯ[�P������o���w�w�}�'̻����x�T��\KtҌ/	4f�ed�����}�|�J�2LnEa���L� �Y�5]#�	�ՐP����Fϫ
;i�j�X�x��9G��Q�9	�L�ț�d�*h��t�
x��Wc����M`:r�]`�q�d�*����s�E2��w�f���gG,hvf���(x�V��<W�-WR�0�	�t�4a)�q��6�H�n������ ����616j���"4R��#���S�[d�k�{��F38�PU��r���FC/���o����*���*�/����/Od�&FGܸ�lB��ǣ~����R]L�}d%$^.�zFӉEw��c�LWA�9��O��i���u�俓���g��w_K&��f��'O��J$�F�����{G�T�56H��,V�F�b��WgM�p�FK2NX�[�c��9
F��5��bi�9�N���N;�;uo^��}�U��ӛ7��ҒC���Si����nZ��)���q�lQg����d�"m �}RG�����%HW�t����)���h X!�w��Y����w�{�[u�>1��yN�\N�f��	I��E�0Y�k���bt�{��Ȃ�m�&k1��C�K^n�#��*6�֙�.���Wj� yh�r��*��H�2F��N)��j�s�	�|�d	�TK0l� I3S��OM�O�J�r`כ�d�"�Lw,�N%$^���+
�eA�Ef��y)5=өE��!x���[�,�g	�}B� <JW�M�[m��"�]�2��_��yEGb����v�zf`�8���	�Y���"hV�����joE��ȼ�U(�b���p��ɹR��-�7&F�&��!i��WÐ�J��P�^��7K�ع̣�$�mbŒA���r�	����î�#��`W�G���	?LZ�G[�2�<�:>{���X"~e����[t���ӂV��H<��գq1�ľS���}��B]DAN���?9�wDd���2+�9��U�{�e��Z�t�F�k�gb`�o���&d^-�2y�������Ϫ�I�ޛd���5b���7_�W+�he'Bz'��W\U-�ld%�v^Ub��Y�l�Ub㳽�ɯt<T�� ����MG=#�7Z�w=ʏ֭�̷���d��i+I�"-�������
lj'��C����v��˕g�;b�������_L�?���y�.�w�Qcb��m`:��a���&��5"لƤ2�hO�ؖ��>����57�'
�}g��{���-$�ϼ>btt�xI���n{]��OE_Q��e+R[BU�,��؂Ԫj�z�,:r���
L��n��1�6$�3�#�od���91ܧ��>����9:�xj�`~?H���S�������!B�NғQ���s��@;7��wnf�?��$�5t+�G�3&`���`�J����=��ܻ�{(�܃R�Չ���Z|R�ټ^�������Z<�� -h�hk^2@�ȼZ��Bn�����c�j��p���,�Ubma|K��������KyD�s���}r���C�Y��<!��QM�#6���<p�6�{I Ə�5��P�B�4����֜��o���h,a�M@+��g���K����B�3_��8�}A؂�,8\0�{:"�~��heݣ�t�z��R��{ C�����GV�]���B�b���o���Fo{D��ĕW�� �e��ˮ]׏�c��9��^ם4Hx@L��tK�#�Hl�W��n-��G�yσ��ZvZ�<�pߨR�7�'ݿ�o�����?�b ��7��8;+�+,7��A�rА�C�3���[����[y��%����W�l��א4�4�B�9}�� ����ɑ�؛5e�>8�v���h/���������=��3P��1ʳH]|�����z������H�$xN�������T�$��`f��Z��j�'�=$SՈ����L'j��ӞA��t�{Ǻi4A�Ě���9��݄:�p�ܨ��^o��V��҆���CRov���&0g�41������X?�q�ǩs)��iS����/����3#���:g�!��J���Hi�Ęs�䨗c�${)''����lU\�����A��J���O��8�%��-d�K�c�b���뺯��p�3>����b^�G���L]\6����☆kB�*��y���,�71U��7��I�d0��^��=L����j�G�Kø��o~�/?c�)�����0����~T���?���z�n�Cv�3�q���\�&�&�L������Gڇ;q�'g�o`!pfi��7J�K�C=&�n|��c����|wzJV�S-�-�u{g�mj����#�HCZ�1�Z6�&0�����W �ž���"���2&��һ��}�ν����>U�vo����L��/�^.�� yw�[�_G��1�4�ǧ'vW��]��od?�T3큅J�о��A����!��t��;z�ny�۔a�<���R�,��m!�[�I@�o�M(ih�@{�������^q��_+V*�:��ٍ:P
"�y<�~-�4rE��˒�}����'���o^Zz���g,_�w����&.��W�&`Iω&%R���[��ڴx�_T��o�]v~�Ĭ�Yh��ժ�M�"@X�9/�7�t^�V��;�����@m�z��4�:8�$��%9?�������Z����2���캶F�T��T�鎣"/������*����;C��4���(d�td电���}%6�W�t�J^�@_�%E�_"��M-5H2~��h?����#�����������ު�Tו?ae��#�9!�������tE�w��RW�˹�SAp�3j3P�� ~fOa_ą]т?il?)��H����a�C�X��G��Bttr�Y�:�"@X<�Qb��؃���4VV�{�����5�#�L�0P䈕(ϻTy�K='���d|�TOA��c���1c�^� �`���;c���V��-��'�^a�)G{@\@6D��J�-�?HϦ�p��k�T�}�'��Y�ې�����U�g�zk����G����N������e����v�������+?|L��t�`;_��ח���궩+����.�72(H
�a��Fk�D�Vz �T����O��ʙ�5t�]w�K��f�2�n�=�*Z�	�,P��x�y2o�Ƭ�P�&��BZ��1����C�x��22��4�X6���V�nߪ�"R�k��
3����I+31��~��u�Wv�A���W�MGЫQ��0u�HA�~Xt����*��o���!Vd��Ԁ��͏��A�(�� �{����V���gSل�	߽�t����z#��|����ĤE�2�y5�_��w�1k��������I�����wy�o���҂������Ape���>�����1�� �l%�t����Z4�<LV=uE�qG��'/�nf��Ҽ �E]+�Oy�z��2�&�Ƹ��1I��}Y�al�-b�ľT}��A�$Cy�F\SG$`��đ��u��W��s��Ťې{�z�W���3���ؘ�l�6�W�nP��@o�C� ��m~�w$��e��f}?��$��}<�y��d��]����Ã�B0��JΎ¾�s%�{�Ek��a��C�b�ŝg��C"�e�|L9�<����j�T|�|��@���E�"n�;E��l�չ#��Bfo3��D��]i���5c����J�a���b���5cm�̒�@�T���k�f��^�3�\P���̬���U� :��F��6Hk��V�!KA�2JP���9=UЫ��O���w����	�Z�P���x63$]�i/(�[�w�ޞ��d{B�7��"x�<$_�L{g�_o��?���?%�4��5I� ��>=6��6*�cC��e��٬S��\��	���]��4�@P�,'�:$ٴIG�M��l�����p<a�*�42��b߄N�6V�E���I��t38K��3��M&)SLY#�/�C����W_�5i�˓�0�(�U����
��l�S��V[�Y���}\�q_�G�C�[+�!
{\V��g��C�${�4������t��%	���֍�.�fCl�����lFO)�tHh��J\�B$=�#i�?��%���_EM���_\wۢ�[�#�;�����h�k?.!�2���w����ޭR���{�_*��>��l�謲	H���7�YG+�c�W�'e���V�~��J��	��s��Y�5�=.���F{+l�}T���!w���(Ѻ�FQ�o��8;�I�k{c2Dxvx��5����u
�%���c�q�8����PA��t>7��翪�᥅�.$4n`�Q�u/Ģ�j^]r��K0]��t�S��v4H6.ʢN��ʮN��[���q�
cE�Tc�,�'�sψ���\���h�{8��%�?����y�~��	A�7��{�}$�9�a�P�����C�t=�[�94蓣�@��W^Ǵ�]46]|-qs�R�*_{H��:���D䈮s$+�m�! y�Ehk��ϲ3�qCe���5r�X�K��X��=���l��v�A��MW��d����`��ա�0y\��~4[d�������릦̶Au��L7�Z=<���O������>8q;g��;ڑܱ��,(D/|�Z4�M�\�<�3*��/�]�L�F_��:�R�5�v��	�I)������S,�&�d��H����{�0�Y���+�꘰�d��Q:��&�*�z�?���1+�1*ZQJ��}1��L��uP�AsZlti
p2�e����0H<pab�cr�Q`�X0�2���MJ�
d����V�0�`�x��u#�bٝk^d��?ľ�N̻�^�t[�m��"6,�%a��#c�4������wT�o)]!��G�]OAị�c%G�
�V�u�5�jO
A'1�y�����"7��=��P���>��wt�3�y�f���@��.m��a�d���m-��6���6(�W�c�.H�AX��na���XY#m��� �U�LW��tB�lU��V�8�^�-��k�^������o�xro���$���6��64��Yg��u��;�W�w�}�Wo��w��f���F��1��kV�۬�%7���!Ɔ�.������5YN3K>�S
x�lE�+�)En�9�ʀ�{ �iYD�9;?�k�z�5��tb:��R�@d��Xh��Z�:�!"Cf�ǌ��߱�X�q}>l泇aŘ�V�ng��Rot����C�א��Wz%��O��?L^�(�OŢ#��Nz6�¤ze���RkG�ĵ`�h(�+j��8����[
�U�О{�Z|ށ�v���OP��=+Y1a�l��¾+b�
����6��AVO�o��M3|�t0�=��!���N&dbhD�P���V*���4��D���Bu%���.�_s|>f��gv�7�lp4o<R(�A9��Z`P"-3��"���Wnf�d��V�3��
�U�[�2X��o���5H(���ֳ�|	�����Ӈ=c@Q�5�J��� ����ƕ�n��tW��.��S����_�M���e}k��m��	�N�F1�w�\��.ϒ)Âg�?	���Wb��ٽ��dT֬�)��Y�/���i�a�V\�M^���n�`�)2J������9B�K#ؕ�d��/��Q5U�A7��V�ag� �"�!����x[�We�Y�BU_ M�5H0�B�+��>�U�z����+��]zx�z͞g[�xC��=n���t]L���z�.��;� �� �5��|')^���>�&ļZy<�_�c��7�H�I���(���v�y�w��x���l/����-���23}��X7O�ߙ ����}��_DK���	���D�g�Z�{��F$� 1l���������	���Y�, Jt0*v���VfƖr�HX�+k�x+�I]�:+��{��(I�[��Cڧf�u�$`��!.X: �c%�$��Dݰ]�\�lڲGK�#΄�G+�1�;���c�i�L����r�e��j0]|u�A��S�Q���*6H�;���觚0�ߙ5Ҁ`'G��<IXw_���ī^^<v�|��`��~	��B`�T�H���V�2)s��VB�o�Кa�Kb����l���˪�����������@��cޠy՗��Z�>�Td���)��#RCm�"�J������ _zfݜ{,f]��Y�J7��][$���&�*����e$�.+=N�k��^-�2$ҷ�?�]�Q���t�=*���We��u�A����o?�KB��ݩ<^?�����{��Nh�������g�"�(�1�(���V�T��������QR��`)��O4)xnJ�9����P��. }i�w&��V7B��zIL؋�����``Y��k�.B�^Q���o�0��׋��t����{�h�J�7s��� ��Z�uF�^W�U`:u���彂�7cV�H#
�nl��^�Q+&�z��䦫�u�Abl��1�}�Nl<yB��\�$�7����!	���Ύ��i�"�sX5������Y�;R��s��7=�]�&V_�����pe���@��8�K� C��W�}#��0s\F�k������h�Q��D�YH�T O�B|$P}/�7��7���p�>���蚗$�g0J_|�7A[� �!��Tg0�'�DSn:)�V�g�:6ݼ`:���t�ƺS����Yr���-�+�,��#a�r߅	�˂g�=�|��;%�-|G{
d'X�̲((�\s��!�E�Ej�H��lՒ-�Y@����t�����۾Ѷ2�{<tx�!�_���c���������g�H�o���=��/�N�(��yS��vո]�F����R`�=�� y��7H�k��#P)�U+R�E�q�*$���
�J�bӍ�L7~�.>~�����f����__n��cQĵǴ#�xq�;[7k�t���s�u	����;h�� Z�;*��	�ݙ���?�R�Y����䰥��w�d�������u�j�~�h�Ñ`�GMI7e\5�Ø>.g��US�s��k����KK���K&ka��D���-J$�{_c�R����D�����s��@$�J��e��t�+��3F��^�p�Q���%$ԑ�i���.���\�_�0���ƢTlه�#��r�Z2W���|�;���wd�}�=I�;�����]��]9��Au�hS����-��y���}PK�$َ�s(JLG����5���`��;�ڪ��Kރ�I��&ǔ�\q9�"g_QRY�E�Y���P�b��(���k(��4�p�>��ʰ>�H	��Vx����[�nY��Q�l���Gde$��T�LeU>6k�2FH�k+�'�D^=�N,�)�tC��W`��R�����c�n���gEj���Ny����'��HH7t�֚��λ���}19*��w�+�]��]\ʚ�m��%ĥ�7`��Ȟ�&�4o$�G��B�����V) ��V��4I��DgT�mLD�"4��r|� Yj�OV�A�"�(f�4Ws3[!�t?�d\x���^jZZ?����C��Np	G�mv��)x�d��� �����J	���t��v�A��1~�֍���$���$������e�2���Нg�Y�\ݿ�R�c=���k �#�X���� psd��&��������d���L��
�od���ض������"���7��83���w��VH����/��f�>�t@��#z_���[��$�>,x�nXpA�>&�q0]|C� �O�İbj8Փu"��J�=�N	t߾�<����Wx���"�w�$�?��"��*�o���N��F���#��;2��Ax/�S�+^c�+�A3�2�!1�ȃ� S������|����*�����eOe&��]/��A���sV�D�}���d:{!�:A��B�hҞ�qE���>�J�*%a7��?ϛ�F0����&E,����zDGЫ��_�B6h�u�jE3H�����O�J���¾�����v�V'�6��h���	8�����l��'Z����Q��]>��C�>&浍M��6�:I�TU)�2��fB��x�h|��vbo�O��M{G`;�W�~�!����_�%Y����7#lR�<�����9+Un�����f^c�Rf���|D97ݏ�M�ry�*����rH�0H��0JL�@t���+e��괇ЌVH�D��1	�{�����-���;-y�Ea]r_�)!�� �������3��zڠg&��!�fܥ�?��Jl�[�<�5�2J�j��R#��̌� ��WDi	���,B�}A�t���!����2�B���v�����_�}Qp�%���� ӱALG�+�D�v�J~:u�ݬ~�/ȳi^18�d4ݐ�n�r�e%$H#vՠ�;JHI6���A'U��yH-2H��{���{��x�ʳJB�Z֮�.y�^���Q��ⓔ~%b$ �)弃}7����97�^m�1��B�m�mh�X����r�'�)���P�>��� a��{8IɅI�@3q��U�9ŧ�:uxH���_y�Z�<���d���[�8:;�U�0)��|n:�ӑ�NA�bӑ�.<���t-4�i�A� 3?�=66��:�u�#?]w`����i�e�����"�w�����MA��:�ɺ�S���;���%�Np�FƤ۔��|���S��(ȫ�&h� ��Q��,wB�͕6iR=�Z�"�8�j(�L�o6Vd��2�=
p�U��TFw�M��� �b��Y<������:W�{9��\�ϡZ��T��z�����)�v�V�M���%����+<[��i�b����ݟ�z�x�wZ�{,�q{��=ө�������$9�n
��L3&��ÞQ�EӡO�*�В��*��z��$����/A��"[�r5HTx��t���J�F�sE����ȭ��M�J�ƨ���f�t��O�w�󓻼U����|�w�+���$A#_�!�$9E���ŷy��1LG5\��ۢu������7tL�_�V!�ܻ���/'!��rL�!�l�j�̓��t�`3J��gIskc��)��������~�4A��D��r5H�
z]V�=�$M(J�y���(Lw�����sO�Q��N�EzUj�������t��4�4��r��@�
�w��ؗ���c���-&�`��e����B�S��?3�t�"-Go�����)�$��0J�XV{D$�}(��h�}#��7��u�J�T����R�Tgh�q�4�1�e|���@���2
٪��A��Whݚ8^��)��A��tV��Ҏ(�U0ݷ��w���l�J7�]6H�t�W��������^S��0���8x��ʳ|gН&dj_j ����^���)܄M���t>�Ҝb�%+C�Z̠IT��4�X��"����~�y��$�p�I��������ā,����V#zg]̹�<C�"l䤣|D��t�n�d��Ԍ14)]!���w*_�^���� <���K��_�ٿ�	2��;��%��űL:$���L����0L�u5�t:l��7�GP6�cC����\��x��x��5"��]�$��U#m�w3Hz��<i��/��~����Zn�6z���W��^*����tg�M��)����P��Jn:�t�Z��7J2H�6�k�Y\��@w��N���,�]��;����#��Y�M&�Ώo��m��l���t1�Va�
��tl�3Y�r����ﮌ�.ޡ��ѧx+A���f�.3��!l�CX���D��[n��e}eT[�n��P�
kq/��.�]�C�B���P���!��š�	��Xp���޷�[�e~�G�Lf���}�̙`+}�B�Z�Y���y�IrFՋ&�ǡ��mPW�g��i�u�w+��{�K�_�p����~��#Mi�tC��f5�G�]v���ߺ�#�T5��@cb>m����ǿt��,��š�Y+#\�����$yLӨ���?�Y�J��0k�k�/���*����j(�27�݇A�Y1YN��,_�,��I�V�ql��8v�6�r��j�=��a6�tj��34�^����f��ư�=E��{�#X�#�q�,���{��{6��#��'Z�Cr"d��^��k�eo^je�K��|�����L��ȣA!$:.M@�T�~��=8�3F�ڪ�:9����@���Ƌ|���?3|Bj-2��qx���&Z�U�Ex�+�v�<��E���C�$mu��I^��b%?�P�"b�FV�B'?��P��{�����#��ΠF>���e�.�U�h��))���:��'�d솖�j��$y���{��d�)$P����j�_5N=DJ~��~+�
g	OW��5G=zq��.�hr�na]cWyh�h��Hy{�Y�����_��5�F;(�qj�v���Y����D���S�D*�8j��s��l�@ԙ�@6�X�F�#����L�l<�7:F��w+}�������öI�(�z$x�����������QF)ԫ�)����o���UI�����aų��0'�Ƙ���>���&F�}Ϯ�)8�X�L �mIo���Ep}�w~��$�����K1�%)���t��u�A�n� �41
l�<m���WM�\�y��^���{\��>��ui�g���Fo-�<�mZY�)г��_��r�������_�]�y�"B �����4;�d.�kz��i�]�4`|��Sw�.��WX���a����k
CCKO���j�{,:�W~%ٚki8{���9�Ӯ$֜E�?�3Uƥ�y_��m���H��G.#�2:��l�4�j�t�iF�@��Ϡ��s�q��O�bj�/������ɪ������\,z?�_�kT/���R=U���M1!~N�*�9�mOK0��2��Y/�#���~�|���lcxc�E���T���Z��[�'��տ�&ǿ�s��d�<�sS]�.����^��d&Γ�U�W_p�9��GՍ]�cf;�Z�v	i�a02=t�hݽ26uS���y�X�"��Ձ������vSm��I-����/�BO)����O��i��U��T�6z�gx?�'�o�Vʦ�K]�Y:Bd>��L^L[]*}���8�P���H�̐�ж��Ja3�x񼬌ϵ��O���l"}����?͛���vo͟��|i�Ak���$TnҲ�{g���[A2ٯzU�e�e�Y��W�uc�j��ݬ�(L)'K]ˤ�.��ෞ����:�I,��k�Yd'��8dF�t����������Fu7�QJ���-���*����J'��0(��C W�h�6 '�Q�9�)W��[�Z��I}�	a �p�s%����o�N`��R�~�;㰅�(bI'6 �(�)q欢zg/�q�\gK�@:ܐ�3Ċ��j�M��}�Sw(�CP�rZRƘ;/�>-(����[�g%h|���JT�+�N&Eǫ��G3T��W��@�U-�����qD��&=����;Ё�P���f����|�>F�;E���]�)���ꨜ@00�"��g̝�D�W���0�i�
U�^g��NЉhy��,���bB�L����ؒ5_1 ���LZOWC2���l@��g�������s#5A2���k�w��=�{q��o�ǜ�j�ru4^��R�oDK�,s�يz-m�B,:x9u��g�Ͱ��A�
��8�u��\Rן�����D3I
5`A:o�r&n�yI}�����_k�ڌ�����:�O\��j�f;!���LS%�&�w{T4��kE9�y4��[�JT<.;d�]��ڤ������m1�)��f����9?77&2�@S�9��@ӿf���;���۫�"� ey�7׹�����*�ո�^˒]�Y�"�F4��}L�Q�u(�]��6*ˎa)� �]i��NЪ���ҸƒT~@X]����h-�eQu�5�%
��"��a3Tyqo���(��y4����̂�vH2J��t�d�lZ[�M,�2?��f�+�O=W9
q���C�������j������ �Fי�;Q���	>��S�9����֢�8l�Kk(�'/��r
�:�� �z��0Va]RV�$[a��M�+s��(������@��}�S��aS�#7OXk�;�5����deW��j�570��73-�c�*��k9t���L<~m9!)t�4��Fc�<���|�/�jR+�(y������K�@�� kuȈ֞�G�^�A����A{܅U�i)ܝEP�7"��̆%3b�Ă��|c�)�O�=����/*~i�(�y�Nu�3\il�cW�j⬝ց0�$�c��'�!k�__+&C��j�_;>
��YP�0W�9~@9�P>WV��)YR��8$�+���1�nόK�)���ڄ�x�������z�$"�8����8�9���Rȷ�g����}ɴ�G���A����l��G~}~��m]��i��N�Z��)�g�Zd2�r보��W���O��_Ce�r:<�)j������'�� "d�+�˽�ʧrT���<#��Т��c�Z�(QW�A��.[�G�9�x�.��3XJ�iD�8|�r�~Z��g�q{�Sk�c�m�Lm)�Nb�/�"M�p�����Ȼ�A�L9�'͹|��Ju�BE�.�����U�D=DY�̤a �m.�nX�ю�{��榙O�.2b��y�l��	e�To������Nr��/�?c�0|���)�|b���mT'?���'r�ٕ&3���t����? �8#�)���s���E���f��
nAb��:O�Lꚑ�/���jѹ+`7�����_U��6�z�+1���d�%��_���f�Y6�D=���ߛ�1�X��7��Gm����7>Yv�TqZ�ϲh� ��|��e��v�3���)U��ʹ���^ҺQ|4��"v����|���	sO_����Tl`d��4�]����0Ŭ3����z���!��Q�<��l:���_}��R��SE��8>gB�4�,*��Ef/�ns�n�dx�0���.�@��!M���G�"g+��/qߚ��O�WF`�޹��P[�3���3g����qW+�3sX�WFj+��yw�� ���i�3AvJ���[$&����;��G������8�Hx�",ہ��@2�L�$��y�(��1-����4V/msV��a�գu�o���׀����$���M���ar}�rD� �?�<QT��%����g�ǉ�O��� +�� xw�V=p����|u����?�w��W����F��4<��o����L���H������&r`:M�ϫȜ[�մ���b��6����m	��s�M �ު_m�w���N9�w�%�c�>#�dR�^�la��n�|L�:���p!�8wɟ���:��߯R	]-��%�����Q��Q��%����Y���W��nW�<�'��8��`�fS�D�J8��8�[�	y��CƷLK�t;O��
����O�L���f$&�}�E�Բ�ĭOB�:�o�\�ֹ���t�_�?��w�hxJ�ҥ�=j]�mx�Tkv8�A�x�:��l�q�]*¢<��U�V�Y�	sdR����%z��`���q8��ս��WY~�A���^d�J�C�C�`�/vKb�.���(�ϽtI�
(3�4�b�
.���s����0���3U��i�ku_@��Y&�OS��F�n�����s��V�bBT߷�=�L#8�:O��|��	��t�S�<T�HK5!͋\��+fn.y3�\�	����@��r��[)����6���r{[�UesZ�q�����`_�A�F� ����d�N�����4�8Z�?�(\��9\�q�c�x�N+f��Lj���Y��RU����O�n�%K�/:c�Jv5Ѥf'~�ǝ�����#4��9>z���ӫ�Ӷ��$�~pF����mb��o�`��G57��Zା[Wͧ�=^H��PR�m�"� ��:��Y
���6!�)8��q���jIge'�X���jag��B���uP7��G1F�?��!�l��2ơ�Y��������Y~��
ϕ�ոA�<�>�P~���U'5%&���R#���U�����,�H���V�\sd<R�F(�H�m�F�g���<c��:�dt�s��n1�[��|G��}Mb����g��U7[�#1��\����"*��t�-~Z�#dv'��ׇ�U��������IU7g
7�����~6���3����d�}u�Ul\���>k_�_?)��y��џ�Γ�:w=��Q��@�^κ!��㗫�v9�],\j��?�Վ���&�ӧ17���D������PQi�*i6���Y�
?�'�o
8 18�ab���k�]��r<x��ڣV�\��#��g�w��*r9ςm����ե�t�C�3�kݯ�k:��QwW^÷����������Ϊ�=ys/��䏭�5!t"����$>���@��^�5�޵޾�Jr��<�ѥ�.M?���3|��Sn1���x��vnH,7_��<�:�b6�*D�Z��,ԪM���O�'w�訹zB�s����>!��ð��V�)o8ͱ�ļ�� 4��oSTs��=T|k7I����	:��}����x}�u`I.�1��.��t�l=����)�uU�Ss�$�o �2���nK�_aF��<B�O.O�X���~{?��ެ�����t���ѫ�Og�;3��v��?�nu$Vf��^	.eB^��5e���3���ݍs�RCӂ�O4�$�-�C;�F��!ZJ�>hj_3�v����G������:j���v�J��p?�7��R�!cYG��n�\i��i�z��PR���z
���-�2q���3zf��u������mo���"x�ؠ�֟K��	%U��������}��A�u%o�tF,��=�J�y���-�BČ+��˓�
�����e�^�R_�Ze��XZݻ�]>��#"v_�v\/�X[��Pز�_��V��8Tج$��z�mE�t��{/��'���x��ZE������ꀝ�u@L�O9�˾�$�E�	`-�����O���= 	����l���������Nt�?,�6���v��R
��/��_B��rwD���=���hY&�I� �gK�� �Xq�2��M��K*����f}x�b?��_��0�/�tV9 ��:?+�G:F(�3�te��K�i}]��;]j&�X��e���f��s��"�F�~>�a�´�R�OL�z�T�߲�c~��� �W�q��r��p],�9��
�:�`�����l��[��l�j}�E8N��zZ�	{-c6GH�S3vc�JY.<�w�m6�iK.��Ft����&�a���LP��D�YY�B_p����ͰH��}ѣƾ���P����[��}L����J]8gm/��5�5��d�_��K�)Q������	�7�ɫ�H�O5+�T�|@����(����ig����B���8�H.Upn�+��[.,:����@) W�_��|"�7����u(&-�8#qg^�Y����҉�E��l�ڀKd��[K.�Z-|��Il��E(�VZ،N+���6h�4�.����~m�.���r�usr��5�A]h4܂
�sL,�T���o�p�]�����|"�F y��/��;��� �y?���B
+��J+��~�*���n��P��B4�VKW�2IX�hd=�{���|�=���ؐb�#�e��miQ��'!5Ks��Q;Q����x��;BE�C�d$>w�!17��m�~��wH`�j���l�r���K�f:Z_]X%��Q�����F.��Io�eS��)�ű�J؀4�R���?J��[�����u�^h/}���뱊6&��ޝM������M6�S�;W��<r���p���y<5Fw��'ue�ӅX��_�^AƜq�Ԁ� ]|��������&z�?Ģ�\���R����k�����_�$՟��WʧX�����`:|R$qyk�[\JѸ3�O��d-��;ˠ7�X>����f�v���N�Z8�)�S�xR�����.�OMV��7r�͗j��Fo��\ʔNT�? �j�[x�>�آ�.�����@�Y�g���y��I�#�=Vn���?��l�{�h9����TIP0�:��� ���l7ļ)i+ħ{��u]��C��I�?�xLUL��P������2h�@�� �����u������=XI��/U�]�zg���w��}�!춪������>��㧰�HJ�?ـ�۩Y��l�`�Ѿ|v�\��O鴹��H��`�[�r�lHz`�s\�Vb�z������	�y/9��8�\7��-M+�i�$�nE~1ƷK�:�`��V�,�o���+��K�l��?>)��P����� ���@\�&|ypgQ�s�p�bm��]�9v�}�	�10�Ϧ7
~7	[���B0V���p�������ۏ���^�p�`8�twd��o��?s��'cn�,�y�Nv5�,�Ǿ֯�.-ع�7*a]�8�o�
 ��x����`|!�c{��Jw�S��|~*?�W�&��~�σ�� �m�F���q��د�-�L���?�ѿ%�W�8�|�z�\� [�V ��F���eE���ZB���l�X��sp}�'�a�#�������)YmutX57Y@PTj�~�,:7f�Rj��Z~F扰J�������t�:z�F��N���{�;�LI]��4�N�,���������5.����QY#��'c����+�q�Sz�
m�,��t�~/�q�_�|k0V�d~�����j�Ђ�.�%����o�P�(t�{Cv�-Ƙ�;zB_����Ҍ�ԾD�� �����u��NsK���Ơi.�p"�kLGۡ�x��W}��jN{��0�+V��~ό�"�R�5�$�$ !jh^��Z��B�%\>[h۸ݲ��R@^�G�����������L��fΒ6�b��9	��(�i��
�4�D�E��	`B�]�Q����F�=�x�ynK��Y��w��i���2�2�c��Ga9�Y����h���u���A颿�c���h���x�K~�34zc��	g3��\Y���2ݐ�'K�R	]�j���$��a�����%W����{\lI���׀ͬ�[~ Z�M�����Ė�c�2��zJ.V�N�N�{��/��nw8����)�^��Y��M2�Qd��3qm�$����B����g��l='v+ ��Z�ь���|��>�)����)c���r��H�������k�����M�v�MLӸ,���i�����-�Ɔ_��X!�,���[ӎ��̧��$�x*��ͿI�jͭ���VJ��@��F�an�LdGb���ӮM��d�va�6l,Y�A�|�-4�H��;o����D��`V�K���8�9�v� �Ʋ�E'~p�h�a���Y�%9o3c-���g�yMt2=��bx����u��l�H�M*q��;s^?^��BU5G�w����~����
ߗcX��'���Բ�����R��\��(��+QxmhQ��d��4&�d���~g���u�vݵ��n����kw�ut����/%K�8h~-od�"R�R0�_�o�_�ڳ����뇁�k��ȃSa��؞-}qL��xe���Т9�j!���c�N�~���;���̝�����W"���m�Y$��=;�Rt��)��|<�&���n���~es9[�-jj����WU�����I@���"��5{�s�2��IC�6<<Ϥ�4P|��*S��V@89���-5��e�EJ0W���$��UPL!>}lQ�l����>Z��<q��@P���;yI�0%��W#�����������0��v}��8s�Sw#V�W}���`���0qKN���\y���s�a����^Z=LLŰ-H��X��G�s����]�d�r�\�D���Fc4���T���H�����P���ܫ�j� S�.�����%>�F.�Jl�4u�u-��X҈̥����4�TX�!�=U�0��[�f��`����R��*���Z����Cwnړ��+�=���x4]@O=�|����%��mғz���������K`�����|�Y����6��Ll��;����3�������1�>w�
�����ءtH��ܴ���<��#^�_3J�Q�1*��,�\ߙ�{�K�v�89�i!��F�Zv�;�Ty�O"L�)�p�7�g_5����WdT���j�!G���Z����l@�(+·GY���0�=�0i֡����-�7-��h�@�m_B��g���s`�������۳d�m�$H0�!���)�2��]~,����K]C���R�&1�B��Y 6�`D���?X)��Cj���em�Lm �w���B��AX��d�G�0��7n`�V�w��:D�!j��#$WP�,Zu[~����$S�Z��#2"�@{H11����u��1�>��1ypr���O��L$��s�J�>e�]R�`�udǞN�^���V�G�u��ݿ����?&CL���`ݓC��vVd�ϣ���x�${�®�/�B�eZ�\�{���J��M�H����A���2�D~���%�����p~XS�ED�5���ȁ�K)N]Q���~W��G|�^��Rl,H&�~6��5�����Dr����Җ��ro'W�`�I\J���{�:!A3
���,�x=Q��D��R\�n1����c¹��zO�k+B�.�ىU�Rqbm1�%��N�x)�*0�'�G �d�VN(��ߛ"���c���
�b���I�.���s-�ښ�f���-ha�'"��^�tY(B�M
g~id�Ɂ�FL�g�ͺ2��0�(���_$�?W��0z�6p�wI���!��j���ݖ�9FA�F׿ͼ�G�lC���x�#��*a�%,���ND��� �hR3�=PZR�f<T��
~*�p�Oi�'K��O`s�g�Sl�����%���&B+��M؞�z@�cr������
%�z������ܰͰ���*�QS���T�H�@�h�|k�����<3ш��	N����@m��N�����[���&c��$Lf5Ѱ��0����v4�C�R����͂�Jq<)�U���G���ݰCXi����6x�ؤ��Zn�`^��WvH��0eզk�a��@n�$������M�Q����O��k���g��{I�V��*���4���B�y���D-����H��S�ƙ .gp�8��F���-4��'4�h�JåؚJ�ѸU�Le��D��K�ZTOYu6��d'�JkՍ 0!m�:�3]�<�\��q��N�%z9�UI�rr�%Ւ�y��Cm
ZG�p(��e�jW��˖��Ol|�$�W���.w��1�d%���l1u!(�������ʩ����-�1�L�]�ʌO}�tqC톞\0m��Hʤ%n�5Y�1C��	
�z4ф��S����w�ܒ��eԈ���L%-#1oF��'GKU�b��rpͮϔ�!ˏ��ǀ�P�h�BB���$��U1��H��EZ,wW�9���l'����Z�+r�EZJ�`�ۅ{� .&aχ'nt>'vz
�tuG��=.y��3���2 �'-XX�ڂ�.Z@m�G��׬S��q����a�U`Г5)Vv@�w6��MH�G��gЩ?4*B����b�-����rb[ه�aj�.�/O�pg/�ΉCU�
�l��<�������Ld@s�6�x��Φ^����  ;���lfe���p�Š�-���Ϋ���|����u['N���-` W/h4�E��A�u�[����gtT����Y��g����������4�R=�fr&j�T㉮�L��Qa��[�M-ǟ`����D�c�X�Y�˕�UZV�1Y�G�F5����MrdV��*��`>���3���/:lF ��J�0-|H��_���?wA�]��ґL��p�����������<����Pn��<	L�=L#��br[q~��|Btq�-[[ֹ���>QB�ZmD�]b+1��T���d�Y��U}��rLrb��l��Vsx�6��e6�"
��������Vjw�d[�� p���~�O��v��5-2�
�:��c��?��w!"�v��{s�7�P3�ꋓa����cs<���?0a�39'Z�>n:�<q� %E�_�5.�wt�0�ݸ�!��p��s��-�g��~�<A�E$
3K��*=W[b�6lk?3����9�)��'�ߙ#�%�c�*��1�Ix8:c��f��M��C���!�7�['��xg�@��ܰY%��*u&�t��I��67 �U��u��Ӊ0�)��cWv:/v񶈂x�	S�Sw�(6��Ы����o�<H�xʣ���1����}���z�Kќ����	��_x��?�l^���3_I"ү�̽uB��f��wR?bTn���z��Z��Xqڬ�-��h�6f�@��X�H����~�V���Mm�A�Zy��`B@L~�a+�E�|az���X�(�K���<j�3��gW���W�|��o��N���)����L��S����^
>b���} ��bS���1"��;�'�=�߬�:�E�?���#v�l�wӡ�a�lƴ���z^~�]V�PƘ�Y��C����n��e��P��Bi��_J�y�
�h��BiT_��6�������~������(���<�<��tk��6l�b�dc��#��--���,�h�b��G<g�Mu�$Ns��Պ��r������� ����5����=Avzeh5!"���n#y*f���~�J��|�;�n�K�{�|CԶvo�H!��E���"v����y�a�C��A��\+:6#?���'t����-?�U�4+m��-�-ٔ�v�A��lY��^�4���=!��G%���.���Z�/��"�߹�q}�/�B��(�!�W`K-���=T���g�V��?�i��w`��T��0�� �8�>ࠤ]G��b>�_��䳯�y����#�̀8Y�zR�kj��[�u��2Y � =N(D)y���?�����I}�_�W�$a����Ȟryf�<mad'�
�=�	�R��T�O
�gP-}n��ϭ��n#���4�L�Ra���켠Yp�6f��:�����g��D�o��L��ƽT�9jX]���s�cӍ?i�F n��<�:���rm�KE%��0ҡ��uuo��EX�Z=��U1���5=ܿ�j}��q���N�N�ȶ�4N&��:6��7���=z�5�����	%f8��u�FǦ��kKlp�md�W�����6/Σ�|���B[��6�>�K����Er3y�!������d��w�/��\E���!Nx��g���n'h���i�p(/鮤���.s����ߴ�r10u,�6�3G���n�r�f�o�Ђ%�������ב������R.���B���1���{�L�6�G��S�H}��nuJ�	���ig�"j3B[�cr����qA��˶�9�ː�nc�?V`3�N�����x�+��#�p6�t�g~���4r�l7�*�Ԥ�C�/�h}J}r ђ�;�����efG����i,M�՜u��p���ߧ�lu9Ln����I��{)ʽ�Q:�S��.n�JO��>`�)����� 㑲��N� K-�'s'7���X!a(;������&�%N�W_�rW/u�>.z�5��)|[g�J��v�����β���z�$����lη"E^jT3!�w�^e�_��!�������ZP^Â�VS.R�^����t�����d�N�,lR�=�)Ď#!׵d�<PA;����]}�|����j���M�Ɏ���ʢI]�~��+�F��ʗ��7��B��fd�Y�pG�ܖ�,�q�]~9���A|-���Z%�=d�nn<9�ad�|�	���S�����j�tq����y!��Բ�Dy��Ƚ;gT���J��z��m��P�W��%+��I:'�K,{������}���$jA9��7�J���|�~�QS��CB�8��������{_��>����U�) �Om��CDƳr������>ۥ�6@p%X�;w����6pȶ�V�A�3m��?[.��:
hw�WֺI�U�ȆX��P/}6���(���zxe����YY������e?��.�(� %j�E8�H�m�w�l�uN6&a�S�H�F���я�rQ��kN:���z�"�4P�ڬ[��G[S�x�E�<��IV���\�;ϑ���C��^<����j�P3j�Jݜx=�ԙvqma�=I_ߍ=;7�T�.�y��&�=�����̳�j���e�{�ܸ�����9X���z�h�}�Qr|�h ����$�4\�4T�a�����V���+�/:Z�w�A�a�N� k�R¼��rZKm��Us�Ӿ�,9�U[AQh{�#�Z,�3(���=s��f1��E'ʩ��f�P���V��l6i U��|���y��j�	��Y�7#�A�|�e�'G#G7%-����!�˄�h�O���<�㔟�Q(��3쉸��R���>cݒ_�Q�i�Ñ[vH���v��뉭�gy�:��րd�b1�������\[Ә6/����ָ��ߡ3�͓4ء|���e	�����F_ȏ�ր��ЖtɓxȀ�o���a_pZr\��3� V�;a�9�2�/��
����0�4V���f'P,�kR�����7Ds�]�O�H$��*�t+$�F_M���J�~�Fe�����9Z����YUĞ��!u,��˙�w��x�f��<��H��\�H�uP7�J ��wW�9����U`�{A�f���C�NM�Dav
V�A̎n����ER��>'C3��9�D�Ȫ%5�L0{��&�B���ȹ�S2���H����l���ڊ8�AV |ꥦY�S
/���^+ª����g1T(Xm����8���D���𴇕6G"m�~t�?�3rd���I&M�m�?���C�<�U���U:�.���R��Cd�w��7ӧQ�+
���0$�J�2��?B�0c"c���s��D�:M��}�]K�jF�K���~WGL{��	K���Ret+��d&��*�F~����Fx�q}6*�&�)N���H���)����1Z~�5su�#p1�1� ��S�b�#�a������F�>�������o[(�#��!�ShH�v
H�����Q?���i� ���j����]!TC��iV�ȳ8���*J9�Wr���C�g���h�����];����iT���� G�A��TX'�h,�P}Z
��=������a5�L�xt��6��
�+)���G��?q����o*��t�~=�d���]`� g��������q"!��r����rw9�E���#�������c/7��g~AO-�uL����C��ˑ=��L�(ѻ�R^yz�#�v�Ȓ�%;
����ȹ�����(�7��xp�<4`=򾱆�?˃$MT�?��Tժ���r�n�`3H�P���z=R�j�9?9\�����7P0�����b.�)(��Q0[F���<��꒏����ʱ$�H���'�D���/@�������ێ�����mm!���Eԧx=Dݫ|��{��nK�؏�XrU�z4c#�m!M�-����T{���b*uV7����c�3�֡��p���~5IJ]X�lCH}qz���Y�p�8�\/�k�=O�"x�T�_>���n�#��Ʒ�7e�-V��KP�Fo0w��{���'E�Iuo=<�;�0t���BZ�CP�>��HP��!D��Le}�Q�b�}z�ʢ�;��~�8�Vln�S�{����]B�	>�gK�L���d�C;~0y�s��ʥ�gÒ�;hmc��"Ch~V�!����<�f��T�ƵzL��?��C*lk@���U/�C0&�GI�_�.ܾ���]�h:[�h|j��#y:�׌�W�:�Ok�=��B��`�,*��Q�R�z����S���4 ���܃����Z�4yz����Jei*�O�ʢ��o��?ۗ�".yu��M`"�-���U�?iI�cKQ�z9��W�o{�̩�U�ɇ�$��Vy���������W�����E�irW�#+JK|�sy"�b��	5�SN���w��$�.6ݸ�Y
>�͖"��dRv�񮭗�y����L���'T.���Mn&V�=K<���x��C���"���z>�pW��yx}��b[�ϖ�AG�q�X8'l��v�Ϳ}��U˰�u�}�e�V,(&'� ѽ�~�~�C@(���H?p��ذ���U��������'x^��e%l�Г������7е������x�4��A���#U`a�@{�9b{����Y���7+,ϔ7s�d&"\�O�����y'���#�&Z�%M�7Sͦ>;N���B*���Ll�����%I)����M���ת�����I���E�cG��T�)���1�U�U�������\�5POR�����t���/�_9|T2^����!g�X�R�a�A�$��?��a��y���}Ai��B������T�`�?PK   ���X��(�O  <X  /   images/4b052587-c364-4d0f-a047-e449c1428d33.png�eT\]�6�,���w�n�CpwK��kp<��;��s�s�yޙ����k5���U�䪫z���(/���� �$%)�����{�9���@(7Q�!R���[�@@H~�O�U��G�=y.	L���K%J�P��^̽-";�PK�}�g}P��WKHc��$XXby���J������̈́\��^;-.+�Czۙ��ׂ.�QE��T8	�DbI��W�b�b��H!`����A���2B���ݞiх��p�7z�?�A������B]����Y��a'�����g�`��
bYLR���S7�#�w���H`�R(������D{��)8�1$�"ބ�#]�����A1 cd��)
��[��D.��j�#md�u���?��wTb���$x�R�!w�~�JN��% �q_A�2�����'>�+�k�)r���{�~B���rw�kU��\�Ð�5\����w6����$�W�
2jY���S���\*�����<w����4���2/�3G��=���Fh�e��d��2�#����C���q3=�|�^�O9o\��쳦23�kL�%��D��޶Y��P;����`C}]�˟3C�j��:��J?�kU��M��W{,���)�9 ��<�ru��/�gY�7nZ��!d�Q�۞K\l2lޕ&��:���?�j������c��A��"��Q����|S4��əkH�
�A��&�"�\fM$�vqE��?�������1��m���Y��o��7�_���a~(���D���TQ4�0{"�Q��!�D(}(�9Y�ޣ@��^���V�Q��1͖s*�kDA��mLk�5�_�	s�i��� ���U3TD��>���Ď���?�Z�W=� o��"��p�X��L�s�%B��� ����`�H+���"�r�f�u��ɡ6�]xsx%�ݰ�v�s��ӈ���տ5��hdv�A�;�0���Q�_�%�0I�ChC8�����a��݆�������u����Z��3l����G.���ͽ�	_�u9D=��4Xΰ�ω��e�3n̚Q3C�g1���enPA{����$5ƨ�(���
4� S�3�t�F����%��ݐ��4=,,,",@6*L [4�l���)��=�&��ؚ���6�8v%���UwJ���x9�� �O\^_�`��[Ձɠ	��I_ki�� ���V_|_zL��t�-�h�N_E,c� �*�`���wU8EI��bŒO:�hfY��}*C|�� ���9��IoL0�N����r�G�?ʉ�����
�5���M��U�ƣ�������T=V{j2�4��iO��D<�KR���РV5W�S�-�V�T�S^.ZȽ�D*�`��}<��شP4$�؀����}#D�Ω�����[�E�K[D�SF$�Ra���V�D�sXtx9�M���#�G���ص�cqfo>���9q䗕�я��OdL1O�O�O�����L����XOLNN��N�Lzd)�P�L��e21�}f��3f2,4��b.e�4�g�f-fk4c�ǣ�!dj��J�K!K�K]b	�;��ɇ�m�6��Cg(֞2g1J2I�NFJ�M�O�I�Ln�-��r?�&m�}$�R�ը�\TU[UzZ�v���7���]���.[=��L�:��&�6��_����ϕ��L�
�x�y�K�����9����[�µ�|���4w#S,/%_+O*�&�w�*=����6�ʏ1mCmoG�O��[?��&�6�<F��d,̺MZ?B�G(0$[&�ѽU��?S��;�:w�U��s���69��)���8:h�l�,k߮��3���*�����̼K���������Y�)2a�����W2�ҫI(���0��a��ތ �e�"!ݢ�o�0HRJ"+��f�ts������2$���\�KU�P�/�6�vt���=5y?xE��k�Ԭ�v�Љ	�-�P�Jn>{�iPKS+0dbFc�e��L�q��u�9|�ؿ<���q�~�~���c7b�mGz:r��KCC]>ɟ�=U��K����Dl~i��ojfjӠ�d���S�S6�E�BlQ�Iu�ֲ��1�y��#Y$�J]�g��L���|������V���)浪2w\�j^�7��k��}�Y��4�8�d}�4�SA��V��Njg4ѣwNw��|����TLEt��.o��>�1b�Wj:���ǖ��r��+�[�>�f%c%U�Z��pB:�G����#�E��Ǩǻ�{�Ս��\�f���=�5�AM�'���/r��-]-1-����/�����K�Z�����)�#/q�:������y�0���6�i����u����wqD��4�����������>-�;{�~������n�V��)�m9gI������|����Jl+����t�`��-Yҩ�e���1�1��%��+�P��d�!nw�{�[���EFT�M���$�f���}凼�:5kF	�V�]i�&��ڒF&]�V��ƍ�j�]���e�Ú#��
���F\��U�֣OMyR�A��.�&�-�^'�щ���+O�[^�������W��<�n?u�}��=���(,z���l�;(m) V D��}�x�O\0�4%�͘�Oû�oy4�]O�I��@xR�1z��6[��x_�@gou~3<�Xv��J�e{�j���?$%#�PMP�'�g����vs��c�^x[�������t�X�m�'m|�H(�(_{<�_U����Y�ϐ��O�#ˬ��?O�!��!�kG�Rk�!�>;���
П�B|�1?z�4A>��wnڦG1e%j!���a�aD	���DS
,'A��A@C�B� g��G ��8$ī?�P!���ܗ���_�?��9��	���Ё�kԿ���Y��=��z�&�""%U��MLl�lq���$AX�/H)e����sUMGM9Y#[kc[CW�O��� ��&�D��V6<��$F� �/�I��q��'єS$��7!�``b`"@ ""�7�(���3��'1st�����������`ko�����������B��wp�q4p��q ��"��#j�`do����ֆ������ɑ���1���� W��J�q�g[�_�02301�]�e���<��&V Qsk�f�Vf>�����:S��9����L����j&�"���cG�������ῆ`�X�?ff���|�}&�P'ӛ��\TA8B�Vi���#�!�S�˽�rR�ª������o�Z{O}|�E��[C����qFue���`���!a�ڀ������&SE�%�C����A3FS�8�[��I�׸T������ɽ�)Ӫ����)k�t���C��#�x�'���&�	�*���"�Ѝ�п��$BL}_���NQ��&��� ��,�h�����^�aA!L �yP����I�--�[w���F�����:!!cw(vb�ɠ����ڠb�
�Z�ل�.Q��٪�����8C�'+�EEEU�a\P�w��j�����?�s�d���Ƥ��QSSO���iTdT�$�pF�������a	�z	}蚜���H��;���˲�� }����r�X(���������A�`�۹�b�5>�ѿ���,�$_�yG$�&�lk�� �B�,i��p�@!q���AO3I�n�9BkP�m�׫��!(�w��������I�Dx���ͷ۩�����j��M�f�oc�l]o�d�\�D�:�?��cB�{��yvX=�}�j:0�ú��s��1��~��_��5�om��d&t�/����<[����	����[��&��ބ�\
�����O'���P2)
�ET���@iz��?�!D���~���t��i�����۷��l���r��}'�d�k�\�t������;3�"�<�ʋ/X�,C�ꮇ��q{�z��BN���K\<�p�A��v�N"�}-�H��P2���^}Ҟe�kd|�L��dz���2-ν����E��Dd�=��6���b�x�Dc�+&�q����x;�M�Ʌ�e)�[52L�������"n���N�6��\�
]�R�JT-���SemV�'n�����X>���r'Xt�Dé�(�rt��rY��Qզ��'ľ�-<��{]6�E�Ǌ0�$���PE��5O����z��V�����$� /�L��d~��t����x�{z ����8���J81"VV
�4���pD�k�Ȧ�-��RbX�e��a��G�ef�������I��諣ŝr���"$��D�D ��k��ĉaX[
J���t=�jY:�.g���*�5��E���������p<�����]�|��X�;.��#��FKS����hc�ҋ`�������"=�d��= �;�!]d�~�MP�o���&�[�KVN��8VAc}H�S��:(�_r�����HȣRRh�Q�s)����XIF&���QV��GS��	�5|��`_#�L�(��!���R������"�.�;U��-kū�B�c�k�j�2ya@˿ٴ��'��P ���d�Sg�c��zk
���\�i �2��Ϻԓ��&��Jh�'C�z)`oa�P:�F�5�s�!�P�zF���eF�Z�:L<�+�T���H��Viu�`hp�]	��.���X����n��BƛB�\�~��_�i�+�v��1�VC�Q� ���.S�In>ǕJ!��.8կ�J@�j���N�؟*�F�gK:����ڭ�;D�������O������?nb,�2cך��[�7g�t��%�9�[ԙ��
��Z��gBW�o+q�p��*��_d��i<����r&�+��V��.zw�`�Gg���m����L1%��v��1��(�kD��,~��8�-h?i��b�0iT��؅�r9�-U�����U�+���Pk	���c��,���9D!�D�M<��t��� "c3���_쭤�J6[�aI�.�&����D ��q:�	���\ޑ#�u�75**�$.��1����N�hiO�-gX<jc%�dddb77�ې,�z�{������+��݌�x,��.����RI��6KZkL��r�.���_ӋC�|�I�8���]VO��r����`F.����=�� �'�¡�JL��^hp(���gB���I����d��_������>���'t�On������7����)0L��W��
0rB����7�!�u;��Ή���w����;�lw-.���q����@1f��:Q/����W�
1�c�$}���-;������0��-'��p\v��V��%K�}Ѥ��&��`����}刿�a��?^�}�^i؍O�¤Ui�x��]0v(�'��{�\B-�_Bo�q�(�C�'�u*�A���FKz�s^M'�+�]��M(kl��c3Z��:��[3_.5A��݊���.�/��(�Iݳȥ���4q��]���Cfu=���֥�C��m�/8�㸡�"�}I�Sc ���@��攗����^�+���w|��b��EjX�ê�Es?��v�dnϿ����bQa�[i�pX������t@0�_xּ� ����P)�4��k�X�`P��7� Kn>ܞs�	/�_}L��f��-�:���m��.hɦa�|�M0��IC�Ȩ7����7A�%4�Ug��D�Bľ���9���}��N7�S�u�<�o,Bb��f���Ȋh_}`LX���`b!ڇ($S�"})�P)B����g��o�wx�B�҈q�`��Հmo�@k���L	�U$0q�DH��Z�8�m���W�
�}
����,���`�h���	��/^q'4�2<��l^̱r�P���|��9 �p9bШ�KC�0��(�_!v�Ky(�Դ�GY�������F[<����J���=`���E]\8rZ�M�qh�g1����&���ڟ)K]�A|�!I2)�Ȱ*�佒�W�i�\�qY��o��,��/�ڄ�=��
��ۡ@��E��s;u K ��t��W.@Vx�����m}b��\���D^�b퉎�ɞ�����;�Op��O�,��R22�E�@��a����'�="mP� ik�i7:R��5][J=��ػ�&
���SPЩ��ܥ��٨����-�V���Ӹ�:�K���������%"��H��:���>�����m�+dKka0R���m�>����se�>|�bMw��3�	�	K�:)�)BDXT?�W�K���s˗��Z�K��Zw�o��<"�^/r�J�u)��]��#U^�k��O��?�1�&�����Z�սu:�7�D�\�Z�~�!�_��Đ�4 o���A���%���<��)W��x6�:p�ܴu>*�t���9f�J@��ȉ�Nk"�S����$�����
�����J~�]��<·f�uִ���3�=�==���LNZ�3���wgZp9q�"��&�zw�hmI���	s�c�|ٲ��)̪b����FȖ��ۇ-ݭ�Dk5 ��a93��F9��� R����r>��b�)9~?}ƠV�-��!����~ȥ�zyto2��������eY�+�ٍ{�]𿁒G�;���?��[�4���ŉ��{~z4�ܟ�M=pB@.`����>׭�J�m{a�o���2�j���{L��}Rfbm� \�f���$	����*���C�ש�$Ie'�	�F�w��/��^����ƕq��F��T��� �B�.��;�>������s�
�a ���]��?�V���/e~�~�����#��.����䥋��,���y<�;.����� ^eT5[o>�[}^�[hw
�(_����״��uq�?ݥ���L|ay�
*}W����|��
mE�]qH�A~~�BE]��w5����G㰔�_̘�W�`ҳ�	_,C�n���T�<f�Q��+�!Oڋ2Y)�贫�Û�-x����C��[�q���H��q,��+��i�������W>L�ㇹ�.�Ȍ��J�z�zv�I|kh�� �����AJ*���8[RG�ț��g�,X �6���}��{o��]�จ�p��qF�������bI]/W�p�2���rii<��O�'D������^+fo�j�Ȅ8u�7�qqq�q[�t�j:�j���&���m1@�>�Z��`�b{�E�o+=����Mx��?��}7`�����&�D�}� 嶉�%yܒ�:�Fx_���[8�Ҍ���wX�_E��3�,�D�fJE��a�{���;���ӹ�d�4z�����ŝ��ˊ��I��z�z�J���S�͹�Ȁc&�?��Qq}[+o�K�5��V�	�x
u�i�2�A�l�HĈ�����L�Vsf�3�j^�~˖% �1�k��<�T���]�s 8{?+��=S��	��C�x��yF�g�����#�������3��"z����{�Y_E�����%��p/��~����:0Y.��OO��幫[���0h�X��4��u�V����S��W%�u1ȼ>pf|>0�G�R%m�w��-���{-Ou?q\jV�V���7�$�Ɩ�^������JZ0$+�~��w��E;GHЮ3sM�6���n��k��K�]=ǝ��Et-D+�F�n�G�yzm޺[�5�O����2C�Q���P�� r��	(�Ex�ּ�IԚ��U�yyns ZIqX/��1��& p)p���o�k��gʴv�������_
x}*<�.��PXƈ�������eq>�/��+t����nh��ч��o^p��
��.a��g�v�~~: ��t�?�J��j��W�i7iM��~�Bg���ϓg�O���v�� ��M�$n�.���kx9�i�a�d��M^Q� 0�b]�Z%��t� ��ЬX<A�stBL�8l<��TĪa!��.��ǲE�4*t�;Sy��D�U��r4K','��ތg>�%mͬ�P���������}WΧ�M2{sbG�,���10ȉ��u8YYU;�&yV:!S� �St���YDX$Pw����lp#K؄��s#�3(*�-�5D�V��%^��
��^��w1JX֭)���,q���2l�d����-~�.Z+��b
�ƽ`��O2!�B� ԝ����y;��Nj=U�4�M"2��჉2����w��X�I��gR���w`y��c�e챹���m4�%0��|V��;Z�-�8Z��ς��Ľ4����Z֏k�  NLNn��{e�?E}}�H�"^�VB!%%�\o���D���e�I�B7��	
����NL�`�� wj��c��}��I�,����G $v'EvP����Ld~c�� _�2u"胡��̎,�o_:+U_}�t't����|�K�� F����@[a%�H��Wjd~fGDH@T��K�ͽ%J��v�*4�q(�{���`�k���k|���x�~0_ut@�W8t�>z
_uՄ�R��l!�б	�}�)�GҢK3#Rg��Z����z�=L�4�{~듡 ��4a�c�}$o^�2
���dO����R��!U��Ww��"RB�8/Fm��F�������u�A>�Ԑ�gD��rZ�c/Qt��Z�����3n��<�7���K���j�eN ��d����ooq)7����`��2K5�?p�����$=�fE����H~�M���H�P�9�����ѽ�|��i�����%�2�̨���f��g݈1�^���9��AvARMe�d#[�5��fŉL|��R��Lg���b��Օ>ܗ[����T��5l�\`X��u�v���O-&�P��<lvq� G40��V����})�sc��3�9{���ٻ�Kw:�z�c�P�p_�e�#Y%���$�4�録��X�+�y�A/nm�������puMS��ф~��$ǌ�9Z4-��|'�����_7)�U�~�s�Uۏ�_^�V��0!�mt�g�x�5�#赕arx��	�+z*�6زYI�d��-�.L��^	�1tR>��-=sPw��U�iG���Y�Ϊ���q��ߋ&y��ґfA�Vw۽�W�X�r·���c�t~ �j'PtW�9p��%-�(�Q���8M �96��i[$t���<��>���Me���~l�̵z'z�����:3�Ԩ{Xb2���,lz,@�4�jY�tL��,i����>kCJm�܋�T�t�\e�n1��??��t�
9�r�q������_�Y���z�:�,�/�>'��6=V����zꑿieE���ߎ��D����Q,��p�D kR�Gf^,�L�K�]� �;m����v+te�f��� �E3��Τ�O�<����;����tv�2�y���Wv�Yg��o"BNES�ǆ��O	2;>�;�7�[�z}���XH��FE�R{��Ǧ�q�6�o�g��"���hP��dR��� ,�2zףv���QX�~�PG����n�8B7�%b����6�O��������e��m�im�e5�䭺5R�xj�����yC��Pfۓ􌋭�\�'�:��+��HZ�r��"Ow2Bӯ�T�)�Nh�kw��W̟Q[0�rڌ�>I\6��d�t�r����[���b���n!��T38xt~NF�۹)���&�݁��f�-�<t�����N�y^������u������o�ң�ʅI��rs\YZs�PS%l�=fv(�����nU�O�#A�|�Q���2�,������szTI�
����s2�L�N>,N�1�,�(�����q5Ɏ�t�f��`�J�w�ĬCOVr[�ul� J�����2I]��%�gԨm]P��ӵ]q�0��z:���ޠ�v�C2���9v��j4��ubm��_��G.	�0�E�>�����ma�݁U.w��X�7.�����Y�.P�����į��6���_ׂ@���7�Tba��X���F����`L8.��X=��>����m%�×!�U�����c�q�X_��2�O�d�)�t��o.VH��+l{r�gi�)k���R�2�V�����ˤ��4!Tx�T�V�&�9J�M�����2mqzv���)d>߀�eT'ߡ�=��Nf�X����S�$�v��U�.�UG�g��0N����rp�HhBՙ�vN�:�w�<�L��]y����|;�+w�l6Xg�?����L� �+�	KG��O�NeoQ�ޛ���Z�ώ��~�#�2YME��Ws�����wn;r9��ZnNܞ���j;��k�N}�LC�Y�RC���úYt^І[Wp��v�R�ע���y���C?�}$ #�:g;׎���U�@�kSt�Rf�9�IG}(�f|ϟ &ܑ��_����d�H5V=��4"3�t&u�����b#��F�1�7��]�8�x�^�
,�;Qm����9�q ���Zp�x�ʢ�X�,��e2�t��f�u�.��%��.��Ʉ�����~l�𪎁���O�q�m�w�QFBs����e��6�k�c������NG�I&�0����L~tj���0�@�)h�β�lzs`�'�Ȣ�ȩm�aPfP���o�)�6MI�d�/�ƃ����#Zd0ev�xw{�ɺT�)�W��r�L:�b�0�wa]���J�<M�7f6>�P����v�����$}rf<6�{
�c�ˋ.L��z��)��a�����߂����{�����7�c�;���&� �ʏ��.�{ND,f����[�e�JE��F����.n�]��3�����Or���i>���$�	�b�$2�R?��?�,�d��Tȍj᧯��Vv�� :�;�CӠ(�Y)y2�����"�T���۳�}_��`+h�%uT!�ҿsT����Ԛ�t��z��>�e{$*\�g�svd.l���a�N�A(�/��=T>,.!7�D�f��-I��f�[~�� >����PA.f�5K�?~�u�ů7E�2���	�H4��?mP�}��w�U+�&�8��8���:����HJ[�����{J������ɅϏ���"X���<���U^]��W{��K>6R�2(5�K����,�33ހ�c��!��K�7���x�ߘ� ����*Fd�}�;���Qq��#Q�O&��J�#���.�`�C_ y�k;.|��j���̺��ld�Q��t�����dA��f�צ�W ��|,?�F�~�r�X��ךH���-�z��6W��Eף�'���e�V!��B�l��>-���Ӄf���V�F���RD �'��Lrn;����:(�+V|]jgZ��\�����溳���������Á�c�������^(��a5-�l ZlL�Cr�x�������YөN��!R�	��Ca��ā�W}�ύ�z�@,�rkG��&�p�	�6�Vܖ�{��]��ܳ}[�˿Nv�//��9�Iu],��|=�5h?ŀ�g(��gU�
ޗ���a�T�f�FQ5P��Ii?����=#�h �BC�6�r�Qz.��B IBU���
���+�6���|�
���j��{�q�����1�-��5��S��#� m�4��9:�y2��4��v�U��,ݓ��zN���0�:Q��P�]�M�tϫ�,!�YgyW�:�k�(~�N���`�P��]�y^˯̣�N�m1ȥ_7�{�'����?;�p���T�b���9P��O!>!Ac��e��8���gT���8�E-���h��T�J��f^{��[�"^~Z.>R�]By�+1f�;�R~���DoӲ��{�
�,�WBW
�su�<�~	[ ���~T>4W���cj'!G��)q�i���.Y��Zq��!��t���p�F��<��o!*sޑQF\:�DjՃ���*I���E��{o�⃓�m���n�G�FmK+��)�����p7YZM�r���sP�&xީvk��/���Z1�,*S�7B<9���
U(i�W�+���i(��G2v}&�yp4"C�e��������}����nd����Ĭ����N�R������p�o��2�����b!��t�Z��'�H)7�(�OR�zG���Ô����6V�桸�gc(=|���5��Un`�ыY��kL�[s��������(���(@��o�ቆ�WcI�'f��-f�{��]?�H�o0��/��a��I�����ks�}���'3��4�a�3N�/2��3�K�e_����W�~|2�u�W����P-����"�Ƨ�_���,�{hv��\��1"SBJ���*�2d��v?W���W{?�U�%�Sݕ�I��nl^O�d��s� ��y�羈S�W����'"��?�=�zܝ�;�}�Oj����0���1�K��]�1�h���<;z{^e�C�����:#a���I���u�@�*_It_�z�h2;�Te�]� �
W��
����b\*���Rǚqj#_��c~ͺ�n��:��zG	N5}$��v3Zef3�Tr��4/_j���/���8̣�����ٝ�[��D��z������c1���k���p���K���B=�H� � +N��SD��g8�LV_0dK�[C�,�"�U������R-E�7OШ�'>W_���LL�_s%�z�9B5J��X9�g�����L�e�&ۜ�EJ��Rx,YD���ՍOK3$~�]�Z��p�tp��i�K^��xNL�ކԂJod�3�mvL[fBm.�	��	ҳr~�,X4��==�r|��yd��d�)?�%@�_|?�)Ŕ��TwZ%PSҳp��M(��t��xzS�ߞr]F.��d^'��~G˥_��H��斬p� Pq0i�W��W�-$�SVSC��� '%����
��n�:tG�ZPTQӻI���8��(B����;ġO=�1�@��q*�׷��rL��A�Q%2=;��yl^��I;�^w5̌	=���0��4Ή[,�=B��b��T+�F㑤���ˋ!��k[ {�I�p��̞�P��m��c��S�T�Kl�Y�Q8�Y$x�/C��#%�1��?K�_?>�����T��t��K��L��ġX&�T�v*�t������X��T�<�&�ֆ��rr�l����9��SGa3��I߰i��)5�Q����}�Ȩ��x2ɩRv���b��"F���kT䁾�ׁ o|��4 v�]�����h�vъ�}����Eo�8�U�e�(£+$�yڲ�9�4��2cU8t����7�;`^1�^��s�%F���NM$���ю:�L9n�hh�l�o'�Q.D�����&�A�?O�����գ�fh%���&xV��Ye�26O�d̈́)=~b�H���6��\�ވ���d�m�1��Tq�5��L+.�𾾘R}[f�C�.�y)���1��v�3Ӡ��x�J,`~���7�I�|�**N��J��W�n�3�L-���n��J�\�ٌ�:{����=ў3�ګ�S�F��Q��-6�x����C(a.~2eԔ>},ue⃯ 2�5_c O��ږ��5�V8����������7���yB�a�d�ݩ�.�pDx���nm�GP��_N�p��m�۝M��M�l��p���o�Qd���T
Iϰ5D��BD7f�M���Q^���o��	ӬJ7̫d9�p����/횿�~�0v&��<�SY	݊����yG��Ō��X���p�,j��XᤠF�������{Q�ּ
k�K]8d�*�}uYW8�'���5�mqT9��U���2h�T��( 9<������x�5�t��8���ǎ%p��p�Q��d���Vm<�<'(�# �q3ۖ��,�ؑ�/}0I���6K-a��O��� ��V�E�LI��8;]�<����$k�
��3�Lj{��ώ��K�l�=��t-�gY;�7�u��Ϭg�������w�$��E���f+�R�R��d��Ӄޝ=���/.�;vǚ�j`q<�96��>�_�,��q=ᱺ���ɞ+c4�S�h��e\ұ���h	�(�_�T���EAT�5[����H�/<[��`�Fw�Dmu� ӚG����)G�*ۯ6�)L9X���Qا�*$*ϣ*F:�ዱ�b�={����1�g2sD�Вg�����D�p�jO^GG�Z��:��O2t!M��7������ ���%~:����Cw�ۖ������Vlrh^W��M�u��r��?:�"^���с��y�:���F�ee[]���ꗞ�-dŒ,Kj�-i���n9Kx��I��EQ��_��*\�*�#]����wG����f����UC��FUI%�{�������U>�CU[;���S�Os���熰;�(<LS,piE�k�x��z,[�W{��7���erj�=8�ϭ���#�s2dH�j�7y��=4�D09+�����2!�Qʻ��}��SK� ���>�J�mۯ�U�K����[i��� )�x:���,~\��!;t䦋7�⾇K�mIl�pb9l�t���7Ih���2���ցF��^�A����:d�^��xe2Ä�cV�"H�K���i��3TpDv����L#ڝ<�A~E�՞�t��o[�Q�ܨ��G'z�j֗��Fӊj���4Ɲ,��fS���\�_���j�:�P6*�,�e88޷U2Z0��U9�(.��>�M�V-)�&i�_em{"q��}V��jwR������8)��e]��ϟo��9 CNTt����d��J�	%k�t�d�!����g,���Qk�Q.N�F��F����w�m��cCf}���[X]�G�^��4/���K^f?3�%4ٰ��ߍx�L|e	�c
ݦ���E�`�ǖ'(�=����������yN����a�ͩ�o�j�BE	��8�ɲ�K,|բ��
�^��߾s?�+�0QT���,��;Za)M6�W�_��m�kKr�Z�\�.������$�����R(^��u�V�{g��b��a��t���ʓQ��g���_1��.��2b|�4Ѷ_]݌y�N2_���@n�T��)��<�]׊c��_td�����S[´, �[t��s�@P+>O��P9/�)�2TcD��&�"�\�%�;$ΰֽ�2;ɨ��Dz�x|=N�Y�E���D��8n��?X�	S�	
VY�\n3��\��p���K�u(K��l�5�d����7��|�^|E���C�a�J䎡�0��K�@סIM<�b�Q�{\\=�J|��}��,��u}��/����a�m�V�kV��v<�؀gs���Xe#B��x
]p��Y�F���xn}����U�U��A�]j�F��4���x;�w��1����^*��V��%/�� ���������4�ʖ�tKk$Ch$�P��L�n�1x8!(f
_�Pf�%��8Pp��\�`�P}}� ��/p����H�@�:��#�� ��h���p2@b��������&B�Z M�Ah|b@4�<$܏�(�z%zM�2��E������R@��I0R����}������J���=�~
�B������QP�~�����"+
X�&��$	�'���
���;pa��e�b�N�1�*_��n� �XJ���_�!G�64��S���E! 14�� o':C@�w �,HLآ��7!��R�l�	<E�� 6����E% �b��������_�r�S=?�
��*~B�;&,W�jD1 ��pd�I^S9�ƄwČ^��Jf���ۚ�GK��$��Xg]�v�o����Zl�!������(��;];-�G�S�;K%nhq.�q�G(r���j��2q78�����CMz�p^�D�����kU-�T�q�%�_�n��Y�1q�R J=�-�Zo����,E��WŹD�$��v�J��������P�N��|2�Ÿuo�����Ki�A�y����\��qҋ.&p�x7(E.�͌�)����mz/��a5q܄yy�Ǩ���s�)����l������Ub��Ϡq�Y$��� |=�w�L*t[:@����i�b�c)eJ��r�R���1�wu8H�	���iQ�J��C�~�aL+X����$~(�_����jG�������ALmb���ӄ၁�2�����Ar^�\XkRA:k
�$����nbXٗ5Q����|�Ij�ۢ8)�����veA��t-2�� �&2(��d`čiR����xy!�d�к�k�.����V�>!�Bmal�� AD�?Q��Q ��`MJ%�ו�Qc5Umw�� ��e�nt:�R+X�<���s���]�3w0�r���2�:����t�.B͟��|����d~u�˷5�16|���#�ᴯ�d�,Z;�b�V��`��R����A��>U�v��e���pҼ�2�����~��z�_�^^���tv�y��Z��ùwu "k�{�����<����p4��iz��F�ek*�yD��ø��&�#|(<3�:�L������I��k����\�S��O�eBx.	�-t����Mżyj�[�7��ʜ��|~���D���!���L�!�0��������ڸJ����z�Y�ǅ���T��4o�=t���U9�ʪ�����)���A �{mҡ�=�6�[�=�K?��~zA;�g�5C��9y��M��ul�t�ny@5�Z�`U�(�X��LG���z6J'�ϝ�9U9�������R~}�%�uz�L�~�m��;���o#��������\;��@�e�壂;��^�<dUc9��!zۻ��Wp�!���̱	z�,��#�V�}ؔ���H��#.k�`�@]��l]�J�|+I��c:�
�ߍxD�#�����XM�2�`�_�v�s�_�ᰙE������c�p�������/�z���W(|k�W;����t%FU�E��R$�D���f��Hh
�]i��&-T���&C�"�� =� F�7*p����뼳g�=3k�Nމ�,���mo��U���1g�C�߬�=����e$~I,��l�
^��zD����V��C��lj��WU�B2���	`�Q3�4�j�T<-� F?���T"��Q�d67�6"�J];���+��ja��hf:�hCRͲ�}��I��{��k��DK��<���@<<�7� a���%�_w��ZzT�8PO�@tX��2R<F��S=V}	Q�*��99��4K��E�ڶ&T�z�P����yNc4A�@Yp�88_�����T2K�[(0�Җ~	w�WF�[b��l�4(���J�1r��&h�=:���P�������԰V%ϙ8�����?ߛ��I�u���8��n�j;���'��\Aj,tY����䐮���*��z=��QT<G�ӕ�>�O���c�N}B[���n�Xhy�����%�~u(��0����y�Nv\����"۪���B�����/��^�}���f�7E���'�צ�DZB�2���_\��eG?`
�������DwV(��"�I����K��euy�)$�q�9I�!���	��Ǖ�K�D/�ҽ7,�s.�"�_� D����L��]]]��	e>:�!��ݥ�$�N[����H��p������ԅJ����������[x�!S���pq�s�=�$�z�N���Z������x�2F�pdQ�,<�a���@_��`|�0�)�(��Q�Nk�LiT	E�1�=��4� CQ�>����
���N����s���p1�T�ԓ+n�a�V�TN넔�c'���g�G��+�@ˈ�w\:{\!�c��\nbb������������� ���~�;�<�P,B�Z^|`�2�cALU��Ki�$�Y��YYA"Y��y�n�!6yHY�sYt�1E��O&�D�H����^�wd_��꾮&�>������zF���Q:����gI��5̦��0pR�Ug8S��t_�ѤZ���ئu��7�}�᲻Ê��1sd�Y$�˼�s�&Hh�BKBmѦ�K(Z����o,�>@ �_��
 -@�{���}���ݓ�L������-"�qH�<C/� �_,��
�=��\xp0K�	�>H���U���Ѯr�����}�m'f��nƢ� ��&�:Wa����2ݝ{z��tKv�v��;�e�F���=��SQI�Ŧ�^�C�6��垳��c���/?�h@�j(D�+��0�&�p����*�H���'6=�9˿��7��
��zl,��Z�:��fiM�ny�Nߌ%f���lI݋�5w�@�C
е@;|X���|�[a�`��e�Z O�c�f�0��[W���/|CS$�a�T �E )s3�k��oK~��>8�S���
�ڞ��&��{�ʢ��T֬�>�ҩ�L��j�F(S�˘jѝ9��� ��O�=!ԱL���W:<��:`U����{rP.�坓��	�Io1��7�e2�ۤڨ��<2���R0��]4B��9O]�����Wd�17�G�ܥ$O
�"�j�B������g�ᔸPֽ�Qa��yu�ԔA~�����7H��x3b�'�&�{��ĳ/E�)<cdS�qg�dY�A�|����u�O �������f
&^��O���X
�C
����>�=D�u��c�	��;��O�x~]>�p!�(�CK�9 ؙ����	���Y"%eZ��n5Z�e�_�4Dk�^lzR7E{~1�+�.�q�t�nѨ�s^�+�C�zdi��o��6��Ũ��;e'
n>�x�an���x�?�t7�/K� z7(4�}�H+�3� �\��兹����sC��^���H�=Pm�A�<S��Op���s[�z�_d�+�� ������|���ݘ<r�t��kS�@]G-�z��^ZP��2����(�қ��G���:������C�8���M�fq/b������|,�1k�١Li�=7�u�y/acqA��͜_���2���t�2�:/7[?0��g�	\��<b��,O
Jtb��>r�J�Ķ��Ց��0jvJ7�K�Y�����U����k�)$�᥄F$��1�jۯ���Ʌ%i�{���L���輐�IF)��m�ɽ4ʅ��0L�8,���S������o	l���m�*=���ruޣ��m1З�эH��o@5}�����-���r �8�ø�����uE�9�
]�����2Y�֡8����`�eB�ᦗe&�k�e�9�/ٵ5G���8���5�e�˘��A׍G!8�[��GgZ����㔽�|��u�k��b�Q���qlJ�Y�%IMn��~D�=��^37�����ґڞ~A�fr^d�n���]�R�����Ű�Gt#n$��;�=5�S���AU�Oc't.�)�6P�ZU�H�3�!�R��������a�B9S^�+�a��03j�r�]g���A��Q����mDښY��p�ʈ��:����~��]��N�����wY�Gjs���WI�I�J�ګ<U�� J�M%�/ZFXk����B��d>�4x��@�rk�>A����\x��. ��=Y�1kD:ɘV^v��|�v'�8��6�� U���~�
R�^����[�&P*+�]
�;���6K*^'�~���X�d(H�k>� z�j�^
�II!���'߆~9�Q�=揢O����J����Ut�)?I�յ����B����p�2�0S�����IRr���zyU�{ylhW��^�n��[�����أ렛����Q��(���]B���ԥIfѿK��3,Ԉ>�]�@S�N�Llyh%B/c����r?�"��i��1Qr"N9:;���POƩ����Nn"fe�%����c�1�<䑺|�-m��������Թ�*�QQ�Jo��ٙ�n���Ҧ�Οԉc�v�mB<�YU2%�M8�T�2m}��'m�P�=\}����b�bc�e��5؈,�����W�����S����#�,Ȕhg��x-���I+����bf�@,�f�zI���������5Wqv̔j=)r>��}������ߪrf�+vqc|܏��� ���z�o��.l�\LTN�D�=x�¾�Y�R���|�+�u��;�W�5��O��m�h���}��qY/�_�o,�0Q$�BHc�U�0����A�_(d����k)c��`\)������x����Y�a>)������*��!��P>ksޣ�(�D�b�3�����Ե��d�V���	��������I��J^-4s��yl�v��͠OcA����q�m=����PK   ���X@��)  /   images/53de0982-6112-45ce-8e57-c75f3734d94a.png�{eWM�5��I�� ��w�;�a��]�kpww'@���;�>0�溟?�~��յ�ԪSGj���Qj_�q�(�p�|�@@@"  �`��롭���w�t��熀����1��
W�,��sރ�ch�!��թb���A&��A怳�>���P1��c4�{?�ԗ̈́�p�i�7�o���q��'Tj��7��+ ��x�t��5��@�4ic����}���R�&�%��_�&D�]���]f3�d�Z��4�����H�Dc��K�j���]tЋ���2������o'*�k7}���������vF��*���g�u�ҴR��FR�(��y�J.���{���>u-y)��ȕ̚���7���/��L�B^��Yz�v���~rm�$�=ھx���%����$�p�(�ێ)�b�d����RW��#|t�#ge������&$5O�v}͎��l�<��էa```v:_��(�m�Xd��!�wgKG�}p�9��q��Z����*��Qp�!S��r0���t{�M�����/*��s�OV���1����3�eȃ0 C1�H�1��Z/[,V��c���~h�~��y�o���}��!V0oڦ���\�#�<��n�����E�v4̥]���<@ �!T���x�ف&dlJà�m������b���-�Ɨ��u�(#x��)���Ŗ��7|x�Z�j�S��(u�2hU����Y��W������ݦ���Ԁ@��Ga߾�X�Qm^�{0xy���pg����w�ל���/[��cu<َi+�u"��ʨ���۳��I�#�Uc�&�[������׉������ܱr����X�rAĈw!��/��6I�˻/Ty�O�R�0�,�8*ɽM*�}�վ���?�kV4ʷ�%�Û��1��[��/uzM�g�P��_a�'y�|�1���!�cQ/ے��恑�x���w��0y���#j^�gX��n�DT}ҨL�@�"9�=H�y_`�~/*�W%�L�kH�3DB�5,�W�@?{���<��������ѻ��껀��	��/b[;��W.�܍d~UI�o�/����R��6�P�wWа,����T�^Nw�A�֪�����%����t��'7��Iy�-�r�|��cC>�܁�������k�8TZh%嘙�k�,lV3�U��{��T��}@���旜�4ӏo��g�.��Bv���sfK=s��:����ʷ���L�1����]�j���1� ��6��uj�[~|�eĔE ���^���/�O~�бd��v�z�7s�2��L��xm�$dr~�t��������L��E4O���q�~�k�9�C$�@«��
0*�9�A-p����"���A�ݻ�ޜ��۟�6�[t�s~U��q��x���}Xń��y��m2ß���É���R����[�gb$Q3�AȆb���$l��TDl��4�m���NIͰ$��te��S	�)��>�9�'���B�Ѐ��k���vgCFt-*�P�ط?eg�Y�ny���N~�
�57{zz=���a�	�ãNݧq:.�"G���-D���e��'7u�\aww���jk㷎wuj,8˚3�"�/?*K��:�%�����v�v2�1�bf(1?���4.�I"ɍǬ��^��k�N���ɢ������"�ථ�T01�Ѝ=�ꊟ��:&2��f~��P�O�Lq�?���N���r��`l�e��ܫI8�������)�,����_��K����>J��r�9Ih~yC���)!���5�н}������[����T�'�-�>*0��ʏwLx�� ���8?�|��PK��O)�I/W.�v�x;�0p�R�l˘�)ո|��,���/��'��:,�d��T������u�b��
��%Br���w?���iI��Q_bu���qՑ\�#���#��(a�t��qeg�� z��"H����l�D���b���.�ө�n��\{[A����a	{Iq&��K�vGm��c��q�h9���
j�h]��<)Iw��q�U����դ�倛j��^ ���������\���D���->�ao��'e�讛���K#��L�FPJ�p���/�_"K0v��5���h�	�80�kw��t�y�V�����U���O�Gl��t4�ʱp�ll?%�!7,5:���n�(�6�,:��F�~��%��OVfJ�z����I��P!�����'�A��F�3���촗��p�(�?T�E݅аA�F��snA�
�ϥ�=�̴�#�b�gV�-�g8����;��'*.U{q��  4E�~���N�I'���P�x��A`�*p���C���Kښ�'��O��A�/6���ކ�5�-'_dD�ۦF����Ά�()��]�KLjQ�E�~NMq* @��5���C][���pQO^x�/�-�&y	��� ���e�lYfʷ�iߝ~�k����}�6z�{t����͞ �N�qC��:;1���ަ0��)�U���vi��C�s���W�C��e�C�t�4��zp�X�_��W�����|�C���Y�å��h,q�W>x����q�������Q���Q%|u� �� �!lg]���i:���x��0�2�p��Trchuy����^@�xiy�+�Aa�N��7���]@4F�&�e��Wl��ȶvu��4��J<�_�a�n���^����h�3� V�ɏ�0����f�N���;��iu�K;~���j�۱�
���	�p�9�����Ew�'11���>{�� ����Xi��n�^^���H��3�@� `���п�jYY(��A�tޠ�������S/�:c��a�l�z9�51��ǡ	���.�ɘ23��K��~�h����~<۹��c`��.-0�`�2B��Ť��M MH�c��2�동k=��y��4ع޻Q�S &&�0����f�~�Dp79y���b�2��L<~�/״���Wz\y�-VSYؓ p��y�5�m��(�uq���{��1��c�ɓ��Oԝ��CK� �4�q�j���Jt�ru��e��c�^�Ӗ��󅤋)�����iP�rp��������Ѱ��K��9��L�����l�J��,����@j�z؀�8��)�����:����P�@��Y��+�;���?��1�p�F_�ϟX����s������>s!;�K�.��?&F2[�i&%�,ߧ��AE�o��U���n'8���?.pr|��~��"�9������Be��t�0��Is��^-�����V�k��]�������~�2����ԗ�\���I�p��Ʋ���0�_g���)�t����N��SR��O�A�O���� �A�酵B)o�&	\��ᖨ�q���?CK)f �����}�Tz�������-wfm�J�ʯ��&T{Y3�E�\r����8[�O�����:L\�A��.�
2���N�;&�i�Ut�����s�e���K��C�
B	W����n���~��NM%�����Δ	[��]DG(9��(Hs0|��T��a>����{L�d���H�ю+�S���ʅ�'$X���P��k�ζ�iS6�huI9g�TݓKև�=�w��$�o����''� �;̽��������q������أ��}�GnȨ�D���Eϭ�z$�mv��C�C�e��a.���}�î�d�"��_:|�y�,4gZ�L�1ɺ�z7P,�eT�_��h�Y��;u=�A4u�U��A����8agF��!�@�� ~7[��k!߷Qg����÷�Da?)�%�UZ���=2X��=o�5�r�+�j3y����s�$Ʈ�}��������*9��2�p�[i����~m�(���n�g��Y��v����h�T�ɔibu�3�T=}�"�MZ�:-6m�_�>G����Ↄ1�C�����Wwt�I���i��f	F��P��8��7��!z�Q��Y䖫*K�_)��z�C�r�;j��v�-�%�%�XNi=�a�[����x��Dww�Ϛ�h����Jj���hQZ�;�|����ܭY��f�
=y�ne����ֽ���X&t������.���t�@ � ,�˂�s�}M8Y���!�� �2"��>���
]��b��@�16����iE���fO��Zz��61�Dg\F��,�N@� ��)舞J�����Mm�O}ɟ�C�`�}�!�7���5it �dC�lL�$�I�@0*`Z9��2��`�x���bM�=9��m��:��?���N�X��u����Q����;�#�ï[�~#Hqi�(�O��P�w���w�����"	���W8�@P�&�u�kg���J���;�z3����{'�&.�����zT^����l2�>M����!UG7>�o_�{��r�&w��/6Ey��~��<kB���׻�N�I�p���f
�&u������C�Ǧ�;����U�1�������iDJ$�w���v!sT;K�=Տ{r���Gj�{hN����q$���ͯ��X#)aG��Gy�^��	�4 �C�	�^�X�&1�O�֫����D)�Fg����S�L!G}���ϼ(nq9�2�tR�+��eF���#؉ey>�NR��g��?��tBy�L�}�Or�:\K��t&�,GY?M[q+1�R'S�Μ�4�G�oֶ`���3����|���d�H!E�BΛ	��.������W�ɪ���!}{q?ڃ{�fl�|�J΁���e�8�ސ��ìs}J_n��R��.���ι�7r/쮎}o���=���0��B4	�
κ��ez�Pބ�O+��MMf�һ����I��3��O6����L�?fn&�ٹ�I&�)�z����= �w;zm�)�'��'|�����\���~ݚ��������>�� �=����L�o��ę�r��{�#½�o�wm�?^���]�s-7��0�B�����$���\�D�O�c������&yG˓���43�6Fcq��dUK�:4����Z�X���(��A����wā���#H2��BLΔ� �u~� .N9w������o�^�u2i�x�5�5��w��<ay4�˳HI�/��y��X�׏�II�D,���Hė�>����S�����S�_䬺i_��'a�e׎3��f�֫G	�?Kо0l$�2�4��,���wItN��f��s]w�=ےqh����o��x�@�|Q2CX0��*o(��r_^Q��ֶ����2vf�=�6hu�B�M���U��;=���s���~	��z8�B��sJ��W��w�Db%�������{��2m�ݗK��w���R����&Q,����U�UL^|�Z�$�%���d�GҫwIC���.����~u=2jc-�e-�U"�mo���9����}?�Y5��8�K��~��b��(dk���#&؉�A2+��4�2��&�(p#�u���^b��}Vt=9�M�q;�u�����S4�9X���N�A�ӗ��(x,'�.��r�j���n�\��K�MI�T�W��2�����u��uP�l�����ّl	K���a҄X� Oc%%�Ж3���J�Sd����R��Yp0�0�tXF����0E�Z�T����� ���#-�B-F�܆�?�]�<�K����o�	�$-3</M�_�N�f̊��~�x��)�Q�En��k���?ĥ9�ZY����x����Ìi�{��d�W2O&E��_���'*�N�
6�+<�.R���S�^�G͊o&BT�7���3K�����ݍ�o�0~�0���Vd���48B�Df8����ƾ��Ѻ�ʑ|r~'�"Bm����wK�lN��b�-�37��:�������h:`h�t�2}���;��-�)
6}h5���LY�� ̓^Mj{����6}�:韬�sX��е���'�W�P�g
�l��LI��g"�P<A�9�a#�w�S|��1�H�8@_�����fP��qQB<��6��
��T��I�as��!S�����S#l��}�t������P�a�蔏���un�(-@��{XV�J�@="��u9�f��6]�8c�π�n�1mڒ����d]�^�h��c�M�֤�8�f y��} ��Q	���x�^�;۸���L��ܢ��:f�$/�駭��B��,��/!��g�cۓ7���:	�%~ �J�O?��������X�sG�</W��Š���f"�
�u�t�fC�s�������4�;tڇ	�c���;B�dF��3F��
s�U���o�KE}�|�	=��9�&�Hs��|�C)���	c��*�n^� �S�y6A��/$=�N�1&K��i0�h����ߩQ��L�\�%ޑ�I�u+'���U�U���/�A/3� :Z�AY#C�{��:M%�5�-�2���h`���B���fϩ,�f�K�� Dc���	W�@'B$7i���#�yDh��IoFb�&��_B�����4�� �#�\c�aA.�%��ھn޷��UjU	,C��^��=��EU�($bP��rq�℈�?���BT�Mm�)�Gj�d��z�㦨�OzG��|��U�}�т� �.����������wb���ٙC,ddD$�hQ���q#�� :�9�1=#�Ȑ�X��Ǵűo����B����v�X����S%S��!�g�VrLo9��/��:}s���~�<���j��h�`D=W�g�������|~\��<va���|?�=�ď��٬<
?�vJ���M�C�
%�� �T�h���>�7~�*�į����ȵ�H($�
�Zn���E��v��g[�?Ĥ:¥L{�Af�b%*�����3T������G�i
ߘ�jih���&��xY�O��fB�,	n*�×}��?��V��NeV̛ X�)�S�';*:�2<8B���:&5��їf+�N����=�V���2��/�)~Չo�u�&��N���v�y*�'����&����޽�\}��O��3�ןf]@��o�VA@�<P��]�:P��1W=���k
9�����5�o���~���b��J������qpW^�W����q3D��GX�a
���9����������d�o�S-|�>KU�@/�J�t���������x��
����shu��}�h���_�����|fv��o�M���I�>SD�K��/]�P|w��=�	7U�2��mv���٢�I�D~���z}��	����g̻�a�&zF�#u�F:��Ʀ�<CHJ�����m�{�|Э��Y�f10z��W+��C�]�Qz@R'a��]/	Q�O�����Gv�k�L~�x�Jn��ʻ�[��y���bI��H�lۗ�8)ώFnE�P�U�[cW��q�y�t��S��9�"�
|X��:[��J�������O�4���d�m�7�q\K�,"y�=�T��	C��'��c�J��ʕ$�&���į��#����1#X����p�E�.Mw].�K����1���	@���87�N�'Lw!6�ۀ�5���=�?D	��F�~�	ن�y���<9f[T�	1+�b+8�m�R�JO��Ũµ��Bgw��?�F*�.\��$�x_#���7��;Yn3�j'�����=]&϶��D��ID�x��>k�7�_c |af*PF!@7S�� @��o��]}i��f?�"x4�IwA7�{y���nwȆ�4�> �.Io�&�p���kަӢ�֌2VبXݘM����X qJ������Z��=1���q/g*0{YY����;��d<�/�����_R���*�[��Vݤ�*�ڜ�fS��O�ʲ1�)N�CɎ�'�������5�bc�s��ID�Ή	�N�u�\����7S�kM�"&\��2ԥ�^:�s��b�#�po"�V'-#������Xkz��^>������FR��Ν&��v� Ix7���^�Cf�� �H����|{�	�Ce2&�?��׵��l9�^"~��o7���C���/K��~O�w�&G/��qvm��(�&uv����7{��Y|3n<�#�Ɂ�Kl������v�X���(��{��!0�2qƪ��\�C��D	f�n��_4����Gx���^&���|"�V�-�N�����/1v}ŕ�����oӉk�]Z�4����_��t�}J&��MP�G�h�	�+��4O����Zy��m����[�^�RXi7kz9��\$v��V-�>�_������Λhp(��:;�{9q]sl��wy���x�	q}���EGA��+Sͫ͒D����A�Y��oG��G5T��E�]-��D�ep/CX�H�QY6��0�ة��hK$���J��N�Ã�C��k7���ON@���,2����l�r�����p-�'J�\���9�����a��e.
B5I���â�s����.*����=�K�?��4�f;�:�׀��B��B�aJ����1V�O�)��/�E��Fmcڟ��}��_��t�l�2��.����1��g������6R�������lN2,8�
�]�S�����S�}U�@X��Ɔ�Mve;��a�0
$��P)}��7#.�T��G\��lp]	>����%t.����V���΍%+[J� �D��h�li��z�X�� nw?�x@%�>JY�x��h�VP��l�Sw~Eji��u����|�M�6���j�^�n�JH�ؿ��dbMߋ�̬�����F��U�!�k\��O	˴�͌7T����r&�m10ͬ�:�j�����ז3fU��Ѳ��W����������E HRBt�U�(�}f!�JBN�,km΂L���HVӦxG 8t���h:�A� /ɒODO;���;�zo�;".�G�,W����%�D:�C1C�5Ŀ@������z)�Ɍ�#�2���OR*dҞ:����ıd�b����t�q���c�׏��q�s�{��RQ��+�ж�mi��s	�l!���UͿ�!�
���)�;�;��Y
c�)�PCp��N�G�_�E;Wh�̲e��	���̲f���56�eV%���e1�~숆�գ��[�+�������R��h��R'��F&��	�@��8�P�'H��E��KX��G"rr�[ZHK�G)�c6R2���=n:�HU�@6��{Q�f�aAb���<��װY�O�}Q6�w*���3��#�����I?I�f��>�%&>4��y� ���VrCｰZe�|x���'Wj��i�o8��e���V��2h}���=�)O�Qe�F2�!�45�L�4ՖuVj�a쫓ρ��j�+$���L�����BU�{�^���T�� :��vYI���
-str�gv�B{t,����kk3�hƃ/�I�'�_%߿��j�v�M 3�ѓOM��D�%�͸N�������z�MD��+���z�@�wL�5t2��_~�c�E�7��G>�w'*3\5�kImt��m���~Oq(^�˘��W¤�z��%7���C;�j����p���v��^N7	a�cz��u�o�j���'a�$��%�7����fQE	6c�c��|Π��|��&� LD\������Pu53asE���z�[_�&�W�@i��D�%���Q��kA�_�4m\��T E��3:���ÄGZ	�@E�YdF���-��>?s�Iz��b��m8�#C[�-�{�뢢!t��!���R����g�1�z��E\���Qly��1sF�;/
l2��g�(e����2`�����H�Bl/!� ��ޏ��ǘ����M�c,W�|��8d0+vP�]$B�v"��GO�����+E�a&$���ћ�P:�>K�P2kŖj��0ߘi������L��o��4�Y{y^t�<6:�V��\�{�}9I~@`��;5�W���o���j�9�ѩ�Q��t���]���k��ΐ�M�7�D�_8�<�C%�[<2��� q�J��ڂ'�B&܅1{�h�����pg�-�^�Z�����*bA�ʭ
#>���+��Bn��d�bksx��x�#}\֜q����|m~�:��'U���A�V-���8=�P*���]	��Є{��9p��Ɵ\�m�ی����o����|{x�[�h����k:�h�f6�>߂����j����<�'�(k�p4��V�I+�$���L��K�5ʿ	��J��l4���t:e��<�9�PU6D\�j��m?[nNp��)�7��.��쑙Q ��uA0��H�Lm��P�ݰ`�1�ixʧS���\a�Y� �~����i����.������|�ɜ��V� �tJvLv=rq�EZ�0+�R�b�nE�G��S+o�V��)-��жx'W~�>3�_[�x�����}�}�z~�ʃ�cQ�C¤��-	 �"$��"��5h���K����g�k�e�$Cjk*�XE}�>�~����וVBVk��'UR>�S����r6����8u3�p���FM}�ԟd���d�n�m?vR�ܼ;�?�~!�l�9�������Ti$�	�vp�}�����>�CөP`�^��,��]�&=5h~�O�{G�O����[�$�G�r������:7Rv�����IF^���9%�L�;���l���&�z�0,�Y��-S:�$���f�	9�)X����8_������O����9�O�k�塩\S�m���B�+X�9�ylI0k�����C�1{�^�� ���-4�8[��8�5N���I^J6sA����ʦ����j�QY������硖�k���M�(���_/uu$#]@�>�$�!�!����Ea��=����fw�>H3�94�Q�]!g3v6*݊4������ǥ)����t��T�_�P���6��~�a.���7",�U�K:�|/���βڶ��]�y�}*�?P��*�~_1�y�.�<���%�L=�-���X���>Ҷ��*M=9��P��od����ck%��x}�ȒMP�I�]	��1mS5�Ҧڝ5O�`L�@卬F�
�%�����7+Pۣk��I��,�G{4BI�0�1�֍�.�K��~��h0�4�E���;˺�~�{����,S�Ѵ��i��=���.%��o�˹�A 6��Z펩��Í�ݿ[�q���9�$M��<q侺ň�����+���������=ʐz~Ffu�X�|�?��}o��K�!p0���ur���8�lD��g�T�>�P7�����a�"3d�3{�
g�������J��%�����|�_#��N������f�j�TO��9=+qT�6�#�L��vf?Rk��|��g���qm������O{�֦<���K�ڝ�E������(u��տd�!�ӗ�A�vi�d݇����f���i7��тG��C���eCX0�h݀��A����'^X����'\�eP+�θz��J��A7�K� u����S~�Z4)��p�W6 �����$�+p�c����`&X��8Q�p��w����Ϸ䠊9�6���A�H�ӗ�u�pV���*}���F���x'�ssd�����1c���{�L�z��R"��o?E}pA����򩓲��Cʜ7���*G_���cv��U%[:٣����|��&��y�|����C�w��fv~]��__�F7H0���$��p<^$��E[BM8�NEG^&�ht.�C$�Q���l�uo�޺��`�4iM�w�q�j���cN9w�5u<ǹd'Y:��n�����.�m~�}S�֥���������x5S�-K��y�����5]G�_�R�-��x`P�8�v�(O�>�n�ݣ,T�XQ����w��������� yR"Y�#l5��`_��ݍغ�G!��f߅�jV��+�����ƴЅ�����
����=��޸ �*
Rj:m�z��>�XS���=:��uy��}F (@�ɽ �X}���p�&Ϩ-��a~'��J�'�:�\}NP�U�&ֽ�m6�n9B�����Z��+�V�[�=���:&���H����ʄ����wR--VX'����kT�g/S��*9 ��T�x�r�L�����J����#v�j15l��H��`����07��gQ-!���@}U��#ƽdL�6Ά��
Ȇ5��?�k�2C�r\`q՗]��b�w���t���yb�h�&`�!�+��k0x�í�ϛ���J�{[K�x�(u�J�Q���j�8q��j��@]"���z�8e�i!�#�Y�Y�1[C�u(��| WuFR��}�S�-�ƹ�0���Q���.�6wm[w$��Z��C7FMЙ���o���ZTnSfv�-a��i\7�φ��_�v��i�u,�eV�;�'ᶔ��B�	��s�a��5g����'|����%���2��\1v�Xk��_G��!��a��H�`����*�41`�~�u���cɈ��t<�	�b����a���0�$��e'1ί���e��c���
���fjg�*�c-z���m���ٚ�����a�fV��ߏ埞�7��-�cfN ���ˊ
��C�+��a��Ѧ��#���a:=i���ݦ]�W�ú�{K6����*�%��d���.�7�y3����-�ʸ����G*��N�Ѳ^�����}L�[��
H�9e���"#Z<��
�F9�6�T�B�ix��P�_�3�̪���W�f1[(��O�|�S����|=�$���b��X��٠�f���:{��J�p��j~��,��-ST�z
=C���+��}�?����X��-�H�k�~�}��XD:I��
�q�h��Dj9�+#D��Z83��På��{��K�?@݂�uq���Tȟ<���J9�!l��|�3#́T�T N_����"�4?���i������0���`����1�n�=�����r�(j�!H^�wp�e�<���\����haBxPXFiY%�Sgd�����f�*�ZH��ɩ2����tƩ�*�(RU+q�h��z��h��/�)ݳ�P�c�SPs�H6���i31�~42�x�Of��l\,���\���x}Y��>9=q�ґS��U�.����<jK�l���l1�#�������m̲�����X��u��Ē�)'�Y��G��}�e�����ū�b�3���n��o�\�G�wį�/m^��P0n�ө\��r�(/~�=4,��.�姚�LCn7AHB�٫~�#�y��cl�qt�*����ApCZS��.fe�s�6������{��BO�<ae:6텖S��:��N��.�Z:0�ͣ������o�(O�����'��f�y"��8���M��q�U�<X�^���>�!R��q��<������z�V�2"���s0�_�5E�HJ��ʿ���P�,5O�!��1��X��7Fq��̔$��j3��w� ���k��[
7��<�E�Ӣ��~��x�B
j�y�I�.yIl��}�-ɌNR�?�$�
�����&LC�DfP��R��J���݆�׈O���Ά��/���,[k�R�yEaQ����3[Ҕ�ڪ�B�l%n�k���@�K��fT�
��ٗ5G,H�ߴ�6r4�id�LB�O�[�j.��e>��f{ġ���@�Ñ$����'���䱳�yl�sZY5��s���5����k���7{� �c�Dqn�C'�q���Љ��S+)1�I&�4W����+u�8D���w�ʴ�s4�Dse���;tQω�{!H��$�����n��P\��n�y�m?���Z.�
5���%���+������/�"Q����K�K';�0+�O_���fpm�ֶ蚾C[%X�Fǳ�	��k��p��/ 5���Ge�K�;\�R�+��2)Ʌb�S��&�kS��R��%>Y�'�M������"��gֲ�����j,���<�K�p���Lz?���(�h���p��X���[zeON��B���J���qSZ%�;/SSr�A��RO�>�g%*V�9K!�����,�M���F�� �ね���ѱ০8��r��wa��'g'���km����G\�Z�Y3:��#�Mp��I��)V�f�֨���ˏ6�z�<#Y+�3�=Z U��Wں��-2⺃��>Ur��|֩^n��n'�Io��D%	Nvr���f2᪣�L�!JÞ���7����[����̖�����SL��tGy��i~�Et��TB6��O�Bz�-V*�A��o�Nb#W��J�,�W;�EZ�h�~-��:��
�H9��i|�
��󝾶Lw(a�x��ZG�(.��<� _�;dּ�5<�?C6���[�D~p��ep"P���4\a<�|�E4��CLT�Gz���P����6~)5�^R��4+�{Oc�m!��U@��s��~#���Ygw�Q:{ԄDA�Hǔj��`�l���m�z�T���^������(��y��yo9(^<iJؠ�X�D�H��~3{�Ze�hz�A/��ܬ&�L� �q�} �#j���U�ea����m�~c��J���l�
�R��3U{��a@ej������7��U����~kz�j���vi��&�h胃F��%=��o�ETYB��&F��l.<?�-I3�t�'aV�D�^�$�~ř����闧U�p�$�d}!q>ah�Ă��~t0�jn����#��)��Uqs���B�����	RH�	Z [��������U�;Lq�t#�*��9�#gCp�mX�B��bj�U4��ݏgY��,�}PZ+���OZ�YMh�l�dH���c1�]�tP-����
�jQ JAq8��|��Ҡzc�Gh#��p|����2�b���QI��H���;
W����	[�e���ALK-є��|�L8Aqrp��s岎z�B��5�Q��0�b·��5�X�H��w�~f� �i�p�Y�~�.ஊEH�4�/}�J�hu�[��1��k/o��|�ߊ�d�cf�AcpWq�M��oJJH���t~u(]�ݚ��F:VV����GL����4��f��'�������G(=Wa��?��)7���`{��P��s5b@ɠ�4	�03��+�߁�pߔWH��^�M%A$^9�>�L�o�NEt8A+�=�?1M�}a���V����ϥ���l�'@a�dI#����h!�H?�M�i��Y��Q�m�y��Sx�%պߙ�!�G��0m���ɓ(�B�n:#	ڹG��$γ q+�x�Ɋ[dO
�)�@y�>yS�-8.:�=�W4�k>�f&NWtO`�^�57H6f25E���vi��4���W��Th��� ���eۣ�ub��h��U�7V�7j��kc�{u��M^Ou����p��}�S�t��KSf�`+�5K�F0��G�-��ݴ%q����2�P��I�D�����-��?�i�j��"�lqln/aQr��[���]�d�XL�B�O�H�F��ڽ�ϣI~�<�H�8�q�9w����-pcRފo�5W�����6����y�_������yhiu/�pS�(WQ!�O��hn�@���r�|�U�Vfٛ��!�㵪�R�+_���6E�f"8�i�)bR�w�p��X�rҹ4�؋�t�vDU}����ΆCo��#���X:#9�.�%��7!��W�d�q�Y�5v[&!�/6�a���&�}Me���5��\�a�$�K3�=�Z��K�y|	�x)v��3h
I�k�8[���CY�9�"-��b��ʲ�8�!�[�ed�Ρ?[��m�gAX��Q_2!�2]+�*�^���_61��ΐ����F���c]׽�J0��;ad��n��|43X�����?g�/r��h�?I�tf���X�f��N7�i���:4�շ���T9�Tɝ�l	�%��5�J�@ա2Yg�t�<ԕL��KO��W��|І"Q��[97�b�;V��K��F�]���}9~��-�
E�AЅ8���e`���5�K�5T�-�J
�� ]��wE���d'�X��Y�{L�Ͻ�/��pd��Х7��ofM�$��n7�n��ƒ�P���z���6kjMx�>!�O��G����D�����do�� �����}v�zﺩᩋ	���=�05s�T8��x���T%`������f�P�F���1���i%�˥�9�`\�&�����Y�s����S�l���k�t�����|rZ����$7���"���C ��	�]ωs+5Nf����0�?t�k:�V�@j5��泥������hƄ��m�"ywc������N+�wa�,��6�9c�%��J�Q ��qx�e	�;x5��������HB�	���$��#*����v�յ�?9"M(��DV~��Z������N�^|�k�S�B���Ch�0�'�	����ŕn�dc|��`@����=���p�NkWm���F+ox�l���@����U=�}�Q�7�I<�`2��� ΑI�R�e���L�J���gA�^��-�ˆ4n��O)@Y.���߹�*���?nnl.���,?w{�e9xn�c�#�g2!�����ԇ�p����� ���֊g�n6jg�ݤ�D��w�k����<B�n�w��ۣb�=��K����O^X���+�.�L͗SOYf�j) �"(�����3��_����L>t��aݭ@����_��X��?�Vv��Y� �\r�B=��u��7+_a�\6�Z����oy�{߫��I�r�����{�<��	A^h�ha��,9Nλ�U��̳����m��fx�^].�`kq�{��y�{6��	���4�!��`��nيSe剧� ����|ꩧ�� ��yh����Zy��U�c2���7�?�,Y�D�z��������؈�E���}W�k��rQ�Ni�\���0����faiٿ�[3xӞm<W����v�1Md�̦$b��6Ԧ @������ܢ{d��sn��`�{3���fdS���s�|<�	�,���eB���mA�&)�x.6*aͨh�����Z���7�n	c
@םq��N*��e��?��I������#��r���m��B%��B���=�a^LJ�l �!����ݽ]
���B\�L�=���fM��j�a�[&˫/�B^{����PA��)�����G��C�ۨO��c��>�6���+L�I'��e���Ym���������a޹���y�0  pL&�(�ʠ0���c��]��ʕ��l�/Z�$�d���+�/��dD.�u{�r��%=��q�O��g�cNF���C悈�2��m���0.S�k�<��s+M�j���)`�`�N2V�"�9Y�Ƶ&Ș]0�7������6�8�E�(x�
�;��m��� �� �XS������/lIg��m���e}gW�(J-f�H�`�H�b��@�iZZ͝�/�5����>�Y�H�U�fLozӛ�G?����|\(8�:H��A�� 
a�1΁�q����{�9���uP�9|ͱ�&n3�!���VѶp,�t��Y|��CK�a����I���h#�YP+�y�+����ʍ���ovъ7�&Յp�={�Q�^�8�S
}�R�`q[�V[�y� �nb�?@��o���<�DW�[锉u��D+�� �mj�Ԩ)Ad�\ 2K�K!�j�Ԩ�ٓ�������S��B���jx>�R�pKoP����s][n����砐!S���r��D%��Z&ǘc;�)hf'�E%�S�;+0"���9���)Ӎ��Sk9�N)�ӎ[_c>3 �$��U�Vi�}��>4z0v|��|@���AK��xZ�ZV¬'Xp��M$��Z����Wf�c�!4�
���`�3�`��orB���I� C kD��=��D�Z]0�0AH�:��4%E��9��&S���q�>���Ae��4Z�ʲ����{��[�Fv��l62�X�ڪڭ��S��؅3�5�	�^1�`Xd�7k��[���1���9q���q�ݾ
��ϸ �}n�}U�c���?X}�|l`ι+�"�u�jSxP萑��\�����cxM*9n\�֔ƋB�D���*�V�}�>G���(u��.>$UyAY3߳f��x�L��@�(iM�V�y��k���Jv��M��.�}�z�ɚ�w/��:a�����^˶`�c}2>B%�c��H�A�������<hR�YK���Cca�F���# Ԣ�_e ��&:M^jVdH�	]F�����'�9�	�&7L=������L�Z�ٔ�4�8���2y��j,�}{wjuC<������c�\Ư��76��zfI�C�ɝ��(�x97�;6���q��Ժ����2p������$L�q��]?�мO��.�A���i�3��j�T�sq� 7��bl���3�q�C����z�TɨR0x��n@V�&ok����3g��!FѪX�3\: d�gRz���ף��F�fQ	����Ý��|Í�p쨔a����G`n�t���o� �7T.�4ak���ΑF��e5@�'��H0X,$�KޠT.EL<ה�����ӛYtA�ܰ*� � ��P�Z�|h2�Ajl�ri�R��Ak��1Q�@��}�?]#��
�4�kt��*8��s5�cw�i����� ������OF�Vo�68:��}��Q%V��;wFnBׂ��B�G�w�n �V�{b����.��2=� \�َ߃\��gD	�p=h�(3 !F��Z0xKbk� �lT�G�؏�DH2/�����*3�Y�ZdAֱ�����ڗ��S�k�PR%ݳRƒ���c�*@��芳�����z�5:�pc�0���G,�`����	�*�q�tsj6oh�R����M�h��z47DD��0Ml�FZ�į� D���8��R��@.�!���q=�H͎.�Lʞ��&C��v,۰)ߨ\�ճ�`��i��/2�t�X&<����oW�4炕S]�>��=�c7�t�n>7�]����;2N0�~UPD���
��Z�h�1F�}�_q����~��������8'��abS��x�-��d<\fH0��,@�0���	����������߯y�k���>C�_���� � 0@�l��Z/A��6��BU�޾^�_ 6
����V��,4�?~��(yYM��֏����
E9w��7ܠ�?ʺCQ���
~���댖�Zfx��s�X��`L`���q�����f��v����L��f
_A��R��B��G퐈�������Zh��k�>{����]��ɧVK�*}���Z�@�YlQ�ޫ�G�;�O"+-��.4-)��) Z�T@W��v�8�Mr�>��`=@��&eB	���q�\��K�.�x7(��+�g���!M����`�{隵�ۼy�BfP���KK��up,�{�'��\ (`�x�5e�b��!��KZT�:��"����F��{����u��S�į�_��g�2�W���rkn�"�g̷E���ݣgq������ *JVٲ�����B�yC)g�E8�T�xp��+�d�a׭��v��B��1*M �����#�礹Z�;q 2w�(�M��Z��+�B�ߥ~!��ν��COjUO�=��%��G�n]���f�$5Ϗ�:�7k�'�#�%������_Z�{��H����6͋[eQk����܋-��$޿�����w߭��:9������&����`ʌS0���Ƞ/��zX8�t� ��f�ƅ@n^������,�×���~���Gq,�����gsv��p<~ñ� �|�I٢�O3v��B��(@�U�u��SOJ�-Z�y��ǩ+4O�e�&��0 o�O����[��`�"7�H�����q�� ���`��S
�M�Av5|��r%u܅� #�@�Ƥ�ZRm��=��<���mL�Nm6�|����n��֐�^2�-���������� ���F�]�IYa��H.0B��B7m,%-�e6=��BW@b79j-6�4��z}�[%�;4�@�k~������� � ���C�	\�0?���� ���r���eP��Q?� 7�k�cG��!�tAo��袱L�U��k|�\U$��2o�+�j�{�N�/�F���	_���%t�Kk	h�����0��ZP�h�q�k�`b"������Bak��?��gRҹq!3�B���es��@n"�L��Ԉ�v�b��ohz����ק@�����\��B���6��w�N��]Q]=V`�B�n����_ށcC��9� ���h���
 �#H���g~�_����0��`&8�����Dt��."ąC2�ߏ�i�L}7�׍Q�� ��pqshE0Ǆ�D�ؖ��h}�0O�/QP�s��5�ǔn�1�u(��^`��5Np�:N��3Q �|}�b�� ǂ�(c@&<��ts<��606��/Aᅟ���TF9wno�C�	����΀�3qӻAN,.|�=>mdsp��:l���.�:V����W얖f�,GG��� �y
}eim�&۷�UV�Ug��:�4�7�X&b�� �(�_{0&OA@���,��l���Q�%��5]j�86;|��3�b��,>�8�b�q-�tuv�0b�<|��l:Zp���5>��I���q< ��d�8����?�=��83�)p4���\�ŭT�ZXcO������9{Y�v=���B9�bE]�%-����C�K_��&��Q����z�9@�C_|����q��P�y�_��7���+����omrq� 6}�4��F.$���k��(���M��f����Ѓ!U�[�R�5&j�4�=X2]ʅ�m�e���Z�X��*�Mii$��w!c���3�ʶ�.���w�[�����I.y�7F�}��`�6���\p��Ua�a��
��[�S&������`� O?1�y�d�T�������k}�k�q�x@�L���7D���Xo�jH� ��J�lI��1
$�V��gl �#Z�`�e,�*af}oݺMv��"�]����݃]M�R���e
J�) "���泮C?���T{���\��J�Pֿ���u��O�r����:��?����#C���T~�\<.' ���+������E�z(��ڵO�=��J��\�Y�[���
T�D�K��֠�. ]L��,uiycMsHd��w�� ���|�)2�?h���oFv	�
����;������#D�v�✘&�����*�87�F���:��lὕ����c�7�	��V!MW_}�Z@���q#c���z�*���O�T�&ċ�̃���@ny�������2�I������c��@c?[��{�V�\�x�\|�%�kj�b����Ui��|�H�P�����B?U�NGx���=��c*�+7��E�h���Z�J���*���\S-����~�'���#��-�j���6Lm�I\<�\��bc�*	Q��N^5��Æ-Is>-My�8У�/� �V�`���m���O���>�}AK��A�:܅ձ����/��PD;L���,Y�9���
,;�5`l4�/���'�|R��c�6���~����y�E�
w\��eR�V���$��K$O�m�����b��\Q��н�w�Cq�����d\L�" =�� �YXXn�9 ��3�0��k����.����|�[���Q������/̾��%G��_)�TE B�GU�T�E:���}�,Eb�=,��P{8�󬲩��la78�Y��M֢�2���������9V˼c�����C<(�^\�%f��N�+t(�2���ɠ���'/��n��C#hmn��^q��^li�k�n)4o�0P<�}�4����Ȏ۴�+�}%�fWC<��(��ۆ�]�2e_q^%b$�p���!�l�fq��$����+��@Ҿ�V�,i�(�b�����j�Ę��4��e�Wv#J�>�'Y� D_4QR`~``�`R[��8n�����׍��w6�p0OM�:��A��q5z� 6e.�U�,m����_�B	��Gg6�j6o�$�=�Z�Ο#���&2}�4Y�dQ�L?%��T��L�h j瀝~�{ߋ~�~�!��@/������#Z�T\p�w����)p\���I^6cW������^�sF;���(H���=��@Qjn�*�Y.��1�A����\�W��@AT ��c2�xr�)��+�kk�Ұ.1��vݻX3hԂns���u���e,�>���eR��C�\�Z]WPf�e3[m�\J�+��P�y�3���>ʲk�G��k��FN;����rQ��:tĚ>}�E\��`B_w�uZ��6�x �IiYpBt�d�1���k}�|��u1V�}�g2ZO�%b�� #�����;8��e��k��$�*d� l2�M��%�nj�����K�:JD��&r���w,Ǎ�!��H����(p�(�+������[*J�P��x�jts@ns<#��<�PD����V	�נ["���-�� ���};d�]j�s6�f	޳��y�	ZP�J���E(8� %��#d�z��}l)��ZO�ׁ9����#����R���׀򁜌׾�r��F��۩ �fË�v���5�'g�q��6�w���$�,��Ϳ.��g��d�Ye��^q��r���F[��"۷o���{��Ӻ�ʁv�9��Ur��ʹ|����>�#��b�]�9>Wl�!�/#ӧ��Ν�d���֔kֆ�U�Zj)ؚ'E���i2�Qb�fj�����H��"p\+����S�fi����X\+�����x��P
���j��j����V���g���XC
V5o֕"���	"���ȃ+}��``��`~Gȧk}��4�9V����B��92T�tQ�X�:��/L�4n乂����VY|�rm�R�x�W�\�I���S5��dI7K���h������_��_���B����&�ʤߞ�EZiHXl��񤣳W�|�qy�чuMa.Qtn���SVi>;���<���Rr�D�b��{�?���̀	[�p��y�*-�Ma��r�}��R� K�_�Z@�`�c`����m�������vO �#,5Lm�f=�7����yg�M2w�B�>m���K��κ��ul]r��À�ϩ�9�?�I�]�>lb�3w�2a$��Dl����1��A7���k-���R��V?��ƅ��!_C��HVz�pu\���� �u�� (�6N�r7�}���h�=��w�c=:�>6n�[9�*���g�]��D�j��=e��*֌��ڦʱ�N5V�d����J;kR�γ��E���S�yGa@X���1�p��1c��-�o�p1G�c��Ռ���J�7��=&;w�0����m�7���O?a��.9�3����SČ`Yt�t`�;���h[�dB��x�J�	�	�g�9�x꼱
:�&�+�}�fО1��+{�w�r�u��	?�St1���2W�[���Ѩ��|�fvw�����d��=�չG{���,r4}�ثha�r��c��m�c�	ƅ&:�h0����5p��D0����̰9Yր��A."��&�t3��Aӊ�@�B��tx0��	 ^�&�L
�=Ρn?Ϗ����ʡ�?�!f{��E�!KL@`�
�O�����H#h��$Jh(ˉ��D3
Z���Ǟ���}.��1��P֘@���f�L6L�j�)����K�h)���z��%��,�[�����1A�Cq<}�c�X���Y��D�pЧ7(w˾����m�Q�ɓ��W6��QZ2���+=����+.����Y�Dݍ��)�!.���'jIg뭫C�M�F�L: l�s�����)��z�̝�n&�7Z��P�����}���
�Ǥ��؄��N�5�&tr��sf1���H���0�L�f�I/V ��u� ��0=TJD�K�KA������e�����S2�K�/� ����7���������N8A��N���ʏ�# ������=�I�e�9I��C����o~3��Z|X�lr������k����w�|��%�i�����uP@Q,��}-�u���J�{�U� x=�����X�F(V+���f�K-�ַ�U_�������{J
�����Z���:�%e��������M4_~oo�TM���^������[.X,��:S�S((�z���@�Ρиg�A�HPH\�S�LW�	S)϶jKy%�:��h�6�J�5��.D�{dR�$ٵ��M���Z%69zw��t�x��~�^�E����NYֲ��im�I.m��r���E�R)!���o#��Z! �XOl6�Q�o�� >C\4�0@�.�G�+��:0Y h���+TS���������|�Ҙ6�]���2�pʤ�
�۷�h�}e�+�����w�B����5�gd)
�qpO`T \�)��������5F�s�O�	0B������
��A�J����j��]pġ���d�_��v�/�˥�2o�!�cm��P4?�s`�̜�D�F�+�i�T���s���SU�?.�7˖/���g�8m�Ƿ��-:�_��Wt�1Gl��?�vwȚ'�ŋ�Ȭ��e�_�4���^�3�=�roi��Ï<(�/]a�grdMn޼�Go�3͢��2P��ф3ƎZ��93�6��l�~�L�fi�e5��VnՒE�Ф#���7��C��\D�?�zܐk-mi���'�o�M�ךg(X �{��- �?c�\'1���h7!���nA5$>Aಅ#}���c������������$8�52W\��MX�((x#@��+��2�� 0Pi��#-���&����wn� �k��q����_/pK��ѳ�>��G�"�@�k%!��6r��D:�@J"�@a�u���%+��_���eS����e��Ge�	�$�d�~�(�j�%~�C!¼3~��}׮
���AX������K��	�פ�:��;�aƻ��ת������̄�
%��n6s>$
�:�q0~�q��=p��A�ɕ�If�E��[�[��,��#BX��Q}���m��_�����;�!g��)���m�ҴԴ�=#T����O�T4,�(�,��%}蔟Ua�����C��J��)*:�p(n������}6wN�4vb��2x���، ��]�	�bW��0��i��������<t���w��C����Ѳ�𾨀pL�}���;��#�{�6D.�����8�pq���RPQ���g�\7���<����p2T#�3�M�6���}u�jv���X�3��N�9k��q����[Rf���=���c�v��U]�{h��Gy$Z[ �0���]�7�e�+����	q,V�| N��b��?�y]������Z�{���}��0���o1������f5�b��S9�M[,9
Be��S�<����� �!͙��f�h�A�*�XHnh
�|.�Bɨܶm՘�״��V|iknU���#!�h��Y��|S����3���G�K%V�g�?d.�r|>��*�4�[4�-pr5f�,1=O&��{@.�хK�̏�w�%�(-���Hp��ܠ,����0��ɀ�c�2l�QQ�x�i�1�D.ѺaN��=����C#�K����@ �4N�ux2Z�1�^��a�a_@1*h�W6g��t^�����+�j6����X`�yͫ��y��A���,�����
���w��	�
����
�2u�qъ�eZ�Q���Y�ip9�I+��9s��!<�2�u�憛��?1��PD7 &�����6���=Ř�U��U4@5%��)��}$PuHW_��Ɛ��877]�(I�m5�!x-$
�ǲ�O|���1Y��t����b�5�͒�޽)�z�t#Д�2�`���M.�����9�x�.��ޣ�&q3MyW�e��������Em��Bf��� *�-��
>gv���;&�1a�P@���ǭ��<�D����/>���?W耈v"S#�g���
5�1�C94���*a�J���߾T��7J��Հn�Q�̝ky�����29mʲn��޿�Eo�EF!	�f�z���h�Y�e]��.C�M�k>���=�ܣ�/�ti	`<�Z'ˌYs/i��gsm��t�î����Im�F �x��3T �,��6�����z��?���v����}{�q�d�tvwȹ�](k_xFt���KS�h�d]f�m�$9jANҹ=2g^��d��ps�Իꪫ���D �����N����(&p<nb��&�M�����}��K�Lj��+����V/�@$bf����"�m�X�~4�u�nj�.4�ڸ���.��L.�P]+­�J���&�1^� �fܺ��5;W��o���� �����(���$өU7&�rqc�u9NC) |>�y\F��	��0Ǆ��Ұc^��B���R���9�|Æ��q`�с���d��^[�Y��ß� �$�L�9��0!�hˈ��4)�w�F�v�ؿ���kUY�AY�9>�' �~��� . ���K˖� [�m��[v(P��y��PpSk��O�5O����j��=,��>'�]���R��~0A�>���<����<��cr��UƼ�&}=�̝�H6o�&���/�*2�\�Yc�Z�ȢE��Y�\����{�N,��/~13�.��ԟl
bLH���vh@��~.:5+添d�ֵB�O�u�����tQ�j!�]MS���tv�� ���ʨ�[��M�'s��7�C�k���A.f�ǻ�DfF�h�E�Z_�8�v���d�|>���j����
@WP��Mܪ�'�I���q��߱E�`;�]��q�R�G�%�g�[!�E*���3{��s�z��^:s)�?��ޒ���<u�t	�e��
��ɀ��Lׅ�Ak,��)Dρ����>��ʧ>�)��~����H�s݊ p}�֚�|�lE�tv�ɶ[e���77	�VI{n4�Q���'���3t��ث(���r��R��_S�!.@�M�[o�뮽Fʥ@��Y �k!V�?��J\$U͘1K��XN9m�6�����[�zu���O�G`����Gsh	`��>�� ��!& �VS{��r�@�y���ӹ_U�\�G�v�����d�
4��2|�h�hM��ۀd0��.�k� 2
��e$W@���x\���s�)��!ƙ5\
W�P�PP��w@�_�}��u�D�w�X^�.)

�q�;D(�-�x�P�k��;}���U���:�@72�0g�8��W(<𗷷O�Y��j= �����E�Sr�+��+�`&�X3��в6Ϭ�q##w��._�ׯ�1�5�\�l߾�X�}�}��������z�{߫�$���]:�)|���_����2c�\��.Es�<����#΀�����rs_S���+*��*R�DP=���o�3���!�U=Sv�L
�&!C���.��~_xѥ�?{oe�Y��>{�]c�IwzHw愐�aPX��̹�8� 
.��\NG�\t)2xQ��W�H!!�$9@�H��t:���w՞��{����U{铳���*յ�7��3��ɮ|���A��� ��l� )����[�����1 �!���x��b��w��k<��M7ڵ�^�X �!�.��m=��-��up�+;�R8;&���%l��Ш�w�;x���-��m�52���aOeSfIZ
�Єc�^�ȩ�6ŋELD�DL�	��]�G�2AYeo��@�*u�T���!b�F���k��*Z�&5�Q(c��)s���i�e3�B*u����F��Ԥ��9�R��Ɲ2���'ռRf�k�~r-��2?�f������v�s.�|;c^Fs��9J���9i:�j��y^��C���G��7�ךA��מ�y%�s�yf���J��9��V��V�c繶�����x��h1oذ��M@�*A��_� ��mp�$�~�sx��\?�?kn\)U\�'������>�r���V�6�\u��$�YPD�	A�B���W9ae�4�O|�U��^�:_L�߳I�� K��ˎ��O�Uw�Z �� ���čMQ
l F�{[>��NMuY�)m����("�
����~"��k��Y���MoT-�)������W�kP�y�G��|�jhb\O��y��R�M~�7�c=T25Ʋod��
�@(�c(�bl<���I���¡�Oe`�!a� �&��0~1.�Ȼ� �^x��)�)�nP�}�	s���'1<1/�m�w+�5�)H4_�#�d
�;��(_�y!g��@���wx��pN�A�λ��]av�����	�2�hS��iw	x+���,�76�s�O�B��u��(M�g�p?4a!H�W\�_G��6m,۶�[�λ��3�mb���pѿ���v�|�8�,*��}���
��b��O�?����ߞv�Ev�3��o���i �$p#M�N>S�3bʂy����ӟ��8t�v���O��o��661ލ��s�p]\���z�T�{eh�U���n��׵��J��C����an1��.�A��.˒b=E�������!'B������pec���k^�':hD����P�5�%�=ER .��'�t!|��_��\�/|�δ�u�J =/{@8�t nDm8��Ĉ�׿�-�})���H��`116���B.?)�?��Ow�������b����"��\!"������'?��o}kW�L5+�M���LEH2�d^ٷ�SjӀ��¼0.��QB}���|����Ks�&��<�&�Q�{�~{��;7�fZQvdHs^g���N��K�p�g'�F)H�Յ�Y8#�S ��d����ǆ�ne��h�n �L��?�|�㡞�x�A0_���&��0¼G���ёh����u_�[o��g�$ʜt-�������������:D��<�h�>_Z������i�س�������wo���ZR�zh���V�~a�F��DȦ�T��ɒ��*t�<]h�v�i�>j{�;<;�\` ��o6�G��=�K��@t�Z��7�Ϋ^�*�w���*�A�%*VyOȑ�F�Ď�Di�H&���qe�� e��3�xS���D8D���!��nਬixaF)E�*ڗ{!���Y�� �C��<�@�#y����(�����B��W�W6\){?�a0A$<${"��#80؊~���=E�A�T?��O�{��^+^bh4�94	4��%�u����&�>�\�T��h�t\C�*����&AP&�ά�C�e>髊�@�`����s��΀�?5d����<}�ޙ[�瓋i�����?������v�3.�y��.4�hƌ���Z��f�_tG�۲�ϱw؇w�xR>��}�s͓���P�%�{�� �� ��D���N�CoP��Nx���uVe��$jB5�i^uhI�i����\��o~�C�!<"F��H�z���F�պ�a(�i���6?;e����>RN�P�s��	�-d?�������AܐH���7T#��T`	6>Ă�90�*ϒ������U$Z�	� ����1�)�"���4���B��Y9�"�����
Q�@s?��ϐ�d���B��{�~q�G?�Qυ�Drg��P�����{��!�H��)��!
��9��ClIj�X�]���ų��r�i�ar�9a�`�h*F������u��z��_�-	��2Ϭ�`42�0P�
q���_�����m�Ͽ��?��cR��kVwn"X�f��:�<�X�AVd��\J�� �V�y�~T���ce]�3�XWi�eQ�W='�j4f՛��꙱9���A��d�	O�����R��O\������K��n�9�HNJ6
B�懀�i{SW����������o8����ol
�8
�d8\��9x�"�mi�����7�CL!(%>��!=��#M�BAuVrۈ(wp/s1�:$q"D)�5�ZE�
��D��k<�k���@���* v܏���X_K���a�1	P�;c�Y8@�t�y/����ғ�E�Y5�-�*/2��nC�@�PY2�DK���Nt��%��w40�>c�Bg.y'��0�Y��~�E�+h|��4h^�	L����ݚ=�c i�B��ǟ9r��*�! a���:�C�AY�琺^�h1�s��w��?�A"~�7~�mx0`L��%�F�)�UB{\�����#f����M��'��N�6��I���I�"�r��>O��xD"/I���&U�������~[D�JQ�,�!�mE��J�ǉ|!@v�j���SL�u�!v"�����|�c�C���5%oh�$�8�X�9��Op,��1�*��sH�Ż ���x����,�i]Fb�R5�hD����^������@Ӑ�esк�/��E����|(�KP!��Ar�鏘&���i��^�W~Z�]9�i���
�VQxDI�k��\�c�b��aj�����p=�DJ��h�p%�;��jt��Ԗ��,��)���t"��V7�R��4Qf[*G!�!g�����<���c�a�s�s����5ߩ`#�I��ƽ���L����	O�����_�Q��æ����}`%?�^UL���>Tw�y��*؛^����R沴EO��/mz�p���ik�w\+��7iK����6�s!����Hlh2��2x'x4� |b��$m��8��Gʂ�+H�Z{f��:�`���,-�#y��� ��Wy�@�U�F�T9�0�a�r�4��B�=�R3�m��N0U�15*s/����+*M��҄�H�Q0ϡ��1m��	舾2F�B"%��&,�Q��#/zFz�41d���\l'$G+I]P%�����t�]�fUA`��|م1�O깕/�܈KQ�V�a�SGm<�{ͺӲ~������u�7��.ɽ���ޑ&�%��`��~�<	�Cc�ӂ>��M	�FZ�[�Q*,�?�'in������{��S�L�Üb��Z�Z�Y����\�����,I��z��m��Al�&g�!�gO��A=B�a��*C��(�=i��w|b�_ �0v�[��C��MQ��H�u!L�7��	B
T!�q��v �0R����4 ��3�:����-oY��h��5���g]B�W����p�.A��	��W�
�]�H� <����?�o��R!-b�3`���	�]f��[����L���O^6��Qqi�3��G�G�W��H?�%#��ɟ�I�����Ea_�y@;0,���3704�R�I�)�6k�=r�H�����^���ʠ�}W�����ϼ}�|�~L$K���=�ަɧ�v�yOw?�b88D�+�]f��	wj�s�6��g�䉖2�4��v�g_�m��i�^z���lP;y�}D��AF�?����L���I�-�0�I���I��,����{�����'�r!��C9�9\(���������S���6���0xB�t�E�$�*��?R5s�����+�} �G��!�Ҡ$#��H	�4���:4�s���Ic]�w�����>C����T�{�L��ES��N����n�U�A|r[Mm!*��� "#kߤ�f��@' 1�h�N{ы^�D��q��I��Aȶ³���=�D�1��Þ�d�D+�ko��-��&��{���	�j�����[��@`Ew���<����&�sS���]�ў}��8\p[Y{�,Ac���pX���h�Ae<���$�)�Ms/�w}���|�z�t&����N�2��Z�W&�7"��7������2���#�
j���1K*����q�/����>w�ҍ���f�o����򐧞&�9��呲5���a��ݞ�-�Qbu��d�4����aʁ���W�b+�'��0�Bd��!���NW�p�ͼc V&�:��Ƚ�T���+!�+	i2��M�7i6��& �5/{ُ{��/�K����9��D"f�䨨bދwRn����e<���K;����L���@��y�ޘc4i�t�w7�|��^S�"K�Y�xўpYe� ��V�P�n�&��Ǳ��C��N6��7�4�3� zu(��EQ�S�KEzt&5\�.��pv��m��aۅ1���^j�X"-ƥr�:W4i`��#���8�,� �A�R�u(!�xSc���_�i&E�=����OїZ���Ķ���V-,8,�CN+���?0�v���61J����*����r6[mXeh�#=Z0W��!�O����$:`y~�w�c+��%ɚ�a
@H��4���"�\)8x� �@���K��O���k�%sL ���X��r��; �MP��e��zJJG��i gA�!���`H�e�8;Fd�A�af�*��@3>�x�≫!^&bN41<s�ԯ�q�T�L�H�H�w��6�w@r0!k���f�5<�5��9Zo���-�
�G�O*��N��bVr�;��/ =@¿��!��5�U��Ԑ`���eƤoT͚<r��AraU�G���i�9?7��[�5�Z$���,��&�E6&�����71��Z��KsHQ1�Ԁ�w�N��\�4��Eӄ��Uׁ�MU���׏B��Y�$�b�z0@��B��b�i���F�-�t�fl�+y5k$�����m���?$��Mws�C��P�š�<����Y��Ɔ����Dh	U�H�X�6Ұ\;S��á�� �a�PA&��5�\�/��H�&pp�Va�;��&� =�@�C�\!Ykp��q��t	؂a �cc W�p���
��3n ps�*��H����0R/'EKRO��@����(݅��T:�9H�0 4$�|��(���YW���,�3<�����K��K]�����ye�06�S��-�CVnm���eײ����92� ��w�C�D@��`E�Z���4�V�Z�l4�*�B-V�Z{7��%�C���=)�]�iHJn(�Q���b� }���L{�@/�?��̘����B#]2�I�,$?lj����	��V�d
o�A`+5A� $�B�� �Ky��c���������I/a�h0B�ɓ��Q�j�l���p!��Ea੯�a4�t�Cͼ@�8�B�P1�H�|�DL��%�mAϒ7�pr��J���c�C���5���x�,$y�m��)���˚DF��cj���H�z ��a,<�Ƹa J�3n�@�8���������9t�'�PAY^���L����B���鏌��v!��k��3֒q�n�
?�Z�y��~��{�\�ϐא�ni����\���{�%�w��J%h;���fg�:׫n�o7��ɝ�';\�nS���$Vp�tzv�Ƃ����Z���H���9̛9��ʜ#����#��,F HL�Zڀ�f�����9�Ym0�r��'�+�<j" *l���o�SŽ9Dlt&�Ŕ���i������jZ��e��C��x�V~F>��}7�a���Lu5�yK|c��#H0�?1iw����34H��`��[��uO%��AG�aH��n8�*�1f�_�-e?_�P�KJ����I�$Bļ*���QZר�[,��3��He��3�+Y�=� �\AT�tǵ��+�>�LM{G��$P�lْ��!�K��Bc~�b�\��()]j�e~蟼E$}
����?0�UQ"�0�sn4.�$� �??����ĝۋ�Z�<����-��� �չ@��묭�,���I�d`rp�f݆��ꗿ2{j_� I�!`�8��k9��R4.Bb3ќ��d�Sռ�`���{f�G�ќ�a���[{��:��I��9�I�b�J�g��CF����F��<0��a���`�fa�	 {���������\�ؖ3և�Ƽ�h����?{�f�7H��M�XS�X�-7���D|�FX�E\�R%;l»M��tjD��|�N��N��4ikj�!M4i�b���I����jj��ׄN�����r��@�"�)!@Wq	�%���(��Ɯ�A��T�L=���IS4{R(?\#_��&�K�&C�[���	�2�,ͷ�M*!��6�[g��M�[�k[��0ng���:�����nrJ��sh8F�N!�=���oe��,�FsL��/�˺p���4ڏ�'R�'�'"��aR���h\��	D�'Xyuq+����˳D���W��Ը(i^�&��Y8�dAA��K���z�-h����>6���06�,��Fk�I��(mR�4Y�]<I�������֞�&	P�H�B�V1K_O�C?MN&)[D��P����B���AjH�O�����.��#@�Z�`�(I_k/��ԅ/��Dr"�i!�t�(�X�g���'iB��S��i��ԦEK������(���X��7�nh.��Rv1}���GK���k �Sg�]����:�ߞ�����/LZ����({-_�.�HZ��3����u�x �/�F|y&���H�hz|Ƴ��F�?��/�$ոE�?|MB��v�����9i�8jRW�I_����_���S�/�ik���[�x��a��3��2�B��B��$���.�"�"_�^WO=�	R�߮�g��`v�У�n�X.��P;�G0~�ż�f����Ŋ{3t�����7�I+��+C�6t��_�Մ��`��萪�ZJ�0��'�OR���Ii),�Fh�����Z ��/%������Hת����;D�b�2슩H��~�@�WذRM�=o�j�� &�k��X;�W z)Õ�"Mn���z�W�DsǵbLi��U�?��_���q9+�<�y��(N�K6>6n��l��yf$;�����ؖh���B���~���C��Ԙ�6H�b�i�.�#��g�g�|Ye�䩛}�Q�����~d��ضc�×##�~�/<�<7��ц�GiH�l;�?zj���	����\eC��9j�>b���ȑ�~�l��9g���=�<zȞ���|�6m�h�~֕��#�2	i�+Y)e��$ &�jË��0�"�b��9�d\��6�o>p{x���i}>�w�˹�<(� ���&K�6��8��_(/!N��K������P�T�m�<�f�K���a���n
��H5�� �.Hc�Y?-I�i��R�R�MR�$i��\wS5=u�L��Ik��9�qN��pa�?f#�9���I$<��w'�@Fa>���g��51�T�*¥yW_Rƥ>�{-Ո�YZ�MPRz����ƹ��J�.���K]>�V7�g�1K�;�-����5:uZeO��Yϵ�G�λ�2�Xw���C6;��e!�;^��
�B���L-�e�i�]�����3�58�����k����s\�����l�Ęu5[�9j߹�[v��~�֎#�7�ȁ��/�/�؞qųm�:k���b/��푽�����,��k�z�&��)��6W�q�.�;�l>�4��O���A;��>.��/���E
%/�p��\�����䬽����D�MN� �]�4G���#.g���(ˮ����x(8ԑ=l�tf�ds�{��o�|�0���f��E|�>Ҵ���#�b�"Rq��FUե6O�KR��G�<�h�B�4��u��_�/Ҕ\H$(��K��Yi)Ϡ����������R9+�Mڀ$s��&�$+�O�	6⹂I$aӔb��� ���������jIpW�N�R!���|�[����J����y���H̓a[���{ ��%���>i�cr<y��E۹�L��-�Çp}��8��`�4B]C�Ƙf�u���'Б'l$���h��q.0nn�a_��ce��_��b��3�+��qx!ur�l#˷��笿��s�*��>��O�5���o�T�u�u����!܁H	a�ڴ��i�z���s׹��<W8j�I��,�^�L�">��J��2�;���Zm��mނ�����unԍ�����OHvP��E��q��4�4�Ţ��;%)�9�fg�!w5<E��sK0^1=S^Tb<o+2l����;����Ѓ�
ߖd)"L���EA�~ˀ�7.�"����~� �ȷ|�!�#C�+�I�`=1 =���q�$6�+��1>b��3�m��o^��)����>o�L����5������	�AzG���uAӃ%K�h�i��3�3�^"���=��^O�G�A�/A�<Y��|�#]�N��-�N�f?���m��u�ٵ�Lв��/"���f�Uw�}����|N��p>�v����bXp_R�nX�6��V��x}�ݻ�m۟�tr�o
WG�=���5[Hw@ �ݜ1|�(	S�n��'�	~+sd/,Ե�|�E^.!}�=ca��0E}���u�~/�⣶������)��.�E#�	��I�٧��޷z=z��SY�p��ށ��@<�ʔ �CH�^�c=nsS,Y�А�R"���W� I�J�,���u#*�\?xa�Q
!�������1����<�f5�?aZ�/V2��� ��q�He�Nޖ�] i�g{��Q��w=9y�6�=y|�M����]�S@w\�O��د��hIr��@�8q%ozӛ|O����M���<�|i����q�w�=g�����졠���]�r�ssպ>r0��z���n\>s�9�o�#�|�=Y���'��N?�f��2�r���b����8a���I� X�����{��zo
�0(=�`.:v�d�=��!'`"n2���4�}"ps-�0�`�>�'�=��s��.�;$q|�\��绑�MWg!X4�#�+R�W!"���!�6�5sĿS<Y�3��P�]����w��`�0r��
��DF^?�����(jᤂ�dw�yH�Ja�A�O],ӄmJ�,����0��]��.�=�iH��M N�ϞZ��f�����r'eS2�e�9�	:_�e{��R5סCm|�~�Xs���(�C�I�x)�d�3Ns;�Ȱ��FAc��_��bm)��w�w]��z��9���g���Ja�y?ϣ#Ѱ\,��~᷂�d���*u�M�l&'<��bXu�
~hk8E���;��[�}�1�Ot�_����Q�[Bɯ$�B����`?s��h�	:IS</ۂ;��Ç�ك��t��@�5N�8!aa��!%����	���$���6��A�<Wf��8Q�[���-�Ik(��B�?��9��t�P����w�RE��P�,�ʮ�g�k�sY��V��!���Agh\��܋�QV��TZ��#��
��&�,6#��;�+�:��AG�ĖD0�]m���ޘ"�~i\u�J���hrm:m�6l���-��~܎�[Z�C���Zr.Xs��C?��:�m�v���\�p{b;�Y�Z�Y"�������:�>��KS�$�H@Nx�?��oL=�rcn�ȿv�v�8�-��f;H�%O�q�~ѓ��\�ŒQ��@-<��o��ou��J�KCB������!*¥�tzϲ-||�}�����+��E��|���/G/�����5E�Bx�f	6.��K�5��1�L��eRq���H�8��Ԡ)b+)�)H�g �@�!��I�yF*&���i�J�8�gTq$h���;c�u
xR�0�,���H{~Aw�;�Q�
B���֑����P�{i��5�N����6�.��'"?��/��~p����k����Ş����u�ξ�w<���۴%F���!������Ǻ@q�{o>h���{�j׭�����S�8����v�#!)���I����F��w����"J��+��:� ��D8�f��Co�Tq�=w��u�z�>���G�p�d�+��6�7����x�8:fa8~֯[k���7o���K�F�8V�z1�R �հ �� /��W�7>�r���� @`��$aJcL��]s��@1ȋԽkm��VµsΚ�fPU+8���2��-Rz�W(u7��`����FcG�A^;���.An�nƌZL���%Ė�����3]b+��&��|� �fL�l��́�3?s�����/^�,cQ�p
��{��Fڀ$��(\��U ���F7<+'�b������3`>Ur�4({��}��r�o�]NPx?������-��|�=���yO�V.U\3��)e�UlR��m!J���ƥ6Jҭ���3
sj��?��n}d�|~�W�ӳ UR�Qğ�E���i�mvg�����u�L�>:T.����mf�������W�ǟ��Uts	�|;�XȾl���0[A���^v�Ka���?�G����	�kQ�B�휟�)�oF�8j���~�E@U��<M d+�X�y�>ג�� H�l�~�n\�@4��~�Xx_���ᣨr����v�H�}���E�\�A�07u�٣�"0�b&�#�0>4��۶�w���a"S%������{đ��q�wv�k����`��,�0����������x�5�$E��������geQ�%�#��<ii���)��3`vc�+̃&�/5?�J� ��!M��������@a�	w�v�=D���`�����e�4�ǿ!H�!�[���"R�1�A�|�(v�2�p��}�=7*j/�-�	-���H��@���y�!���:���hI�'�e}��7��6�=�-���z�LO�ځ'{�#y��y��a	
��=��0��[�U��<B>4b+���B���x�A�ǎ�5Q�9g���89;r8�yb|�7.�g�{�My,���@_���F2Z���	۾�b����c��[��={
svȃ6{[��<i#|�U�� _�ڇ�Py�]��gن��mnv��ز�n?x�8=0���䙢��u�]yՋ|s�H,"��� j x0đM�	�x��?di1x�Æ������TPM�?}4�&�B=H9��7!D#��0�:!�kæ�c%�l�����@�k�l��aO$��Ę\-��9�Jf��a`���^Z�$ߴ@����:�%��7}�N ���b�� d;�w�G���CCX$� -�F^Z���y䅣��`�ߺ¯��n	����A+��F)�~C(0C@�
�/�q��ay.̅��YCT�O����uF��؉2YMa�J��ܰU��)b�zr-�C���E����>go�h<�a��/�@�U�����!�̟� ���P�<�g�NU�V׎]�b1��|5��#AZ�gsӁ ����
w�Q�+K��o�F�2B�Π;��+�)�N	A(c��p�Q�,F�<���)[�R�P_������oۺ+KwrȎNO�����OJ��9��߲y����/��Ns�$���vXj9��v��܀���5��l�����e��l��.xz؈�@?�X �U���۶�U�}�o�ѱxp�q�-`�&iR
�#i��?b�㏹��(V`p������!�'�?�CA�ǵ4l�|ۍH�Vؼ�J �@���ߍ, ��-w_��yA���ɼra�b����Z�x��H�lP�~`.儗�(�g��"� ����9$�)I�)���T��I�o�&8���AH���3���'��a�;�d�L��W-����@Z�����u�J&�� �E����7@��?��%Mr��~��k��� ��?����!���3�:0��"Θ ^0�MK�씌�uG�e�L�RV3/�a�d+e@U<wU����|�}����"G�ћ�^w�u��[�Rd���0ƶvݨ5֌�qT���[��� ���5�܂s�p>��͠C�3������y�u&��'��[�/����#�$�}���+���Mm�94g��k��=j��DOd�ư��watj8��h+���w��[Bɓm'<�Ԕ7}��	/�@�<O�����>������7�����U��x�Y�����-��@ H8<O�B��<3��g+��"�Lĵl$
�R:�Z���5ힻo�COl��Բf#fW���G����׾�]�<Z�T�20����Ԅq*~�"z�c	BB2�o�)/D7�Ad��H��F�5N��HT�$E��Y*j!��4Kg
�(��pPyh`���� /��#El*�k��͡
d�J����GՉ����>���9hE������"B$d� ��{�k ����_��B����a�XO�-��3�
�u0vy.)/3~��++�F�f��"L�70���Zs��G� 2����'�����=�;��,���y�� �ӷ˯x��>���֊R�ds�A����6;�̈V�W�U+�%y#{��d�>�����^��Z�����l;���W<�r+W
����gO��2���{l��=���;β��0�s66�ƾ��o���E���&�_��I[�:���Zu�֎G�M^�z�i_��F��Q鐺0����x��Ojz)l�@H<�Z�y���`S(=C��G��`q_n�]�u�ɥdU��k������ᾩ���Q�)�V5F4�[��3|�˓��≯�����UP�M�S�����T�����Vau�9)���)���q�D"T�C��	���i?��-��`R���ai��Ռ?����>�p�yS9l���i���^�g�p{�rL��F�V��)g�4D�[j[`�� %K+Ax���)�.Ps���N�����ξD�C���Ʌ�w ��H(������.���<��"s��!ӟ�Tu-���H�vl9h	��%Z�iI�?��ʖpO�3Ʒ��Q�Wݏ>��(�@8K�h�/�>�-�~#��I��<�e��W����0���w��{~���s��;�|�^b� �0g��@|��p>�v�eW��݀A��@?#���/}���_ז�P�����-�S�ֺ�폎�I���l^6�E]l�u��9;K Ҽcmn$�t\��$k>C��lⷿ����t����jc�[���o ���d�%��qVZ$�`�c65��L!+��-0���{0x��y2�h��-���k�Xz���p�qGc3C�f����Z��	���F�����!L���<@`�/�\�t_�B(���hi}U1gɨ�ajt_v�d>�V�z��`��Щ�������ijo�zB ���M�M\X3c��)����x��|x���<����%h�w �5�ɳ?��O!`���{�����+�3�:ׁ�C�!�h�q��ٻhPt��|�рphh�|�f���rb��>���_�^D�	��D�zZ�|����<p�9d��4�ݤ~���.�S�}C�!!��J���0��/p)��$���������|��a����_���-�ܵ��5�����2`Y�J|p�}#st )h5c�1���������h��:����7?_��x�v?��}�߿�v|d43�M��$��O]���N�����	���#	pPq9�GZ��_x���� y�J�ݖ���_�5,"y����A�}r�3�T6���_�MsU��[�!�܀- 	��i$�N��,��=�q8D^:H�H�ܧ���ڇ/djoJ,i�Xq��P�t�P5�����9������,����RJ����
�������b���]���d��F�	?��s�q/*���9���n�!���ј�Ӂ�	��0�o}�[�>��@�T���@$��e�<���<�Ϙ3�@��<%~|��0����m�>���o���<�,T�JB �g��Ә+�=�va\.�7��wF�^��=" բ<�A=H���Ʒ�F��uߧ}�Z��@P�]F�1v��_�_��~����(@�g�g�D}RT��cM����;�~Ͼ��[��`�w�3�y�B�A�~؞x��� ��'��rWЅ���C�?����QJb�:����&�`�>�s���\�&G�T�M��o��$d�H��ˠ�$��H�HLHe
�`��y(+d7�K�0�з�vچM6;w8�;���Tp[>���+�,y�k���^��(�'_~�����W�jw��N'���d�|���$?�Y�zQ��?�;�`��.UJJ�f���V�y?X5�1��H�iV��I+��@0ހ�0��� �!�z�_�NEf��yF��i Ҵ�r&�њ~\���\p7�̃�} n�� 8,NhG��U^�����}�<,���F̃
��{���T��Y�����_Q�i-
e>�[���
�×�I��{�5i�*��r�`�%A^*���%L]X�ny��9��zιچ����ѽ�������-�:.,�m�M�؍??�`�\���GJ�C�Ё!���M8�gl$�RΆ��8 ��R��F.�^�crk�0�'���}Z��s�V�\I��v⛷�!*`�<�l�NW"���A�'��z���| ³�9{�k_c?��{�U�q5�|!��L��Ar�4��ԋc8vQB�{�"�JC�q۸aKP'��X<&9���k�{)Q��د F�=�2��G�w�t8�O��?��/��s����{�<���v?�ֽ�E��?j\~�3��P�E?�B�^�Cب$0Ta0i���A��N{�e9)4�t�s��t�0�2�ʯ?��&��'���^{�΄xv���(+k~���p~������u׸0	��+Ulnf֦'��?�
������;��soz�y���/{�;��5���R�.����4׿`(E��9�ŰR��bR~����Zנ9CH#������,;m'�B�K]S)Y��|�����sA�:g��߸�=|:n(�sO퉖��6 GyF�0Tj�Ԣ(�Ja���c�q���ȜH{!y�sWo��`��sG:Y_�8��u�s�棞\�n#h�=+)�<�*|'<��*��R�ۖ�< ��7�������"�}�tM"@��#��
��:��Kv�X���Ar��q������"щͥ�h@jogѦ�7M!�R� B���1�~�����ʴ	�La�O����Z�]Z�\�
&�'D���P����*�U�&L����	J�z ��|8���Z�x"��5�,�f@���ۉ�	GNSU�,$z�w\f��q�N���;I�����g�����M� ~r7A>9;�{����TԆ�����B�Q��%,��[��'h��k���b��ҡ�\�RB�+t�#M�j�
ԔP�����۹��.�b��9U�}�������mQZY�EF4{���#������w��!�w`�$UEH䝣w,�:64��
�p���t�q������L���=�W�L�`؃>C� ���z`��4ߗ�+0�Ft,FDy�H2^v~���]�ΡZ+7��g�k"�\�;6����3��#��3������F��)"��n<�u�!aT��S6��
b�Y�<0"�C%gx9D^�00
�h>��3�A��Nޖ�ow��T�b�� �i5�iz"����l|�tX�u�+�=yȓK�&��z�U�.$)�Cl��[,��ڮ~�����+p>	i��5���c��=��l/q��V�'�	_`I�;�x�V��p���\}�cӶb�u��!�$�S��S��I��x$�
�Z���_�B����=�Vn2|��+����O��r0s�T��SЄl$�z��?(& R�ŝ�.>�&����&���G}�:�$L|�B�f������O��HS+MAƋ�ϻa x~!$ +��\|��/�4}�7Z� o��峂E<15C4 �ߵ���m���)%J��R1�0̑�#Vܷ�6���6b#k�ݘ�̗��A������Gr�T!�ԾM�4��*���qg���V|�O���\�rZ�4�*�*q������+xBը�3/�(�5MӪ�J�<�n�������=V��
.�P6[��s80(��
̢m�����ʃ��̻K'�+�B$�~M����J�P�Ӡ���ru��M��V�&�=-+)�1~�S�{h�N*wG(�N~i�"����Q�$d��]i!t���1�g�����!�4 ŀ�]� Oa��y���7�_���o�t���N�Ȗĉ���j��ٓ�r�������u�6�E^�q�}�8B[����p�����mG�J��jZ�+x�����m��I�5�-��޶ԋD��K���t>$]��<$$��`���\"�z�H�0Vmn��~�d'�y9:L�8E�0$r��<_I��X��c-��@�d������=���2p��VjE4��DL!�Z.�YZ��\W���ؽG�f����!u�@�U�K_W���Y�HN���i�g0FEz��k��%�IWM>LHbh��0ϐ�41e,=բg4�Z���px�N���x5k��o�38bs�i/��C	E?�H���`m�s�s�+Pp�m�A���~�	R[M;�u\M<q%�+�E�_���(:+O�]>�*�-���I�4a������?���\ j�	+H�5��0��b;��t�d/��uJ��!��k�@��-��iv	P��ޗ������.3M��p�r$"t҆�Ҽ8+51NͯR�^pt�,��ȴ&����LS�5a��GYYaH$$�xs��"%����"�a�J��E_�R�UeA��Q%2�gb'o�jQݞ���A�G$.,���P{?�z0<�H�{)����T�+0����ƂI "Ÿ�|��Śq}�d���=j�� �!w�=�1��l�_����?7�����vq�*cq8#l�\ڌT�M��$�*Ǐ2=�Z�4F`%�*� -ō�v�el�dÕ��$���F���6�U83ӳAI
?��Ē��V�9%]��%b�������@ɾ!C�r�H�#�m#WB�C��[IЋ<md3P�v�B�Xk&�Hާ<@b ����$�9�v�
`�$e��+6D����������j��N�&AFn��ߒh�Å?<b��~g �5'ؕ�׿.�x����]�/_tXO��D��|�U�����,Ы�A{���D����K���^e��TX�=y��'�9�_�è2*|;����(����cc1hfzzƯ��"
u4���`Iz��O	�
�N�`~f��w/���$��m�}��wY�Q'l�V݉?Iܦ��V��(�V��%��2�����?{|V����� �:�҂䛾��%>�)��Y�J�����vi��
^i��C��u_��O����`���=���Dwzf�/xL�.5"�܄uMZ'���=�Y�s�r%�ڹX�qdl�|U�ȉU4��n��,PP,�S���i6cpY������������Ҧݽ��w$/��^ӑD���y�7�Ʃ@�d�	O�;�)�^��C<U���g�s�:�FFǭ�P�#A�{�὞��۾��݅k��H��+zR��P4)yO�Y�������U¦��29{#��byh�3��N7챃�V]h�T�(��V�+���]iW�טSb�B9��k��Ȩz��jO��ǟ}��J7�,I<�j 6��Mw�P���oqfn��5�]��O��aÒg�`��H�7�C&c�����Od�cCn�y�[~���B�]8�k\�)��'�
���ύ����$���B��֬�Ds3s���cl20����ƀ=i���N�d-�2�	?�Ǘ�>
?;�>�xW��S�n�/��]~�v��A���K�/���4��
]����`�dt�_\�E���na�Hl�tNۢ��i[�U\�y�G�N���U����;<56���1�!5�۱�Ѡ����)��j+����S�O�w��%ҔN-O�'���Y�EϋB���Yg���m۶%�Ջ���!��9'�F'0�3�\:<kÕ	�K��+�3�,�w�K�/�}�C��L�#��!�I���{�� ��fi��3�lu�����);K��k�(4;�o���Z����j����)[����� �/��\��>�����]#l�:���h�T)Lz�"��ٺ��ڦ�6xpɸ���|%���7�t�둵��E��"�*�n�N3t���C�BP]�^l&o��ݲѱ���uWu�T�fe��"�?}ih��(<<M� ����+��jA[��O��o�|��%�L�����\��᜔����yخC�q�����G&�����\��0⮝Ĳ���l
�D��Q i�3M]�r�'�}�G�񩐓\}_��W�}dk-�"�E�!��l�zz`L[����rm$©O~�N|�?��@6D{��?a�#�dW��S;�������q�0p�g=�6>����Nد���{��'WA��{��^_�`7�s�N��_�e�5'E .}^�7�@HS���FU-@�Hi6h%*�%����s �'�-�������0���I�"���*F���T�[s����ک֧-c ���O�<V�˓�$\�-x����CONNۚ��6::�I�<-J�-����b��b������zh��>�������)�&�lg��L��5��}s8�s6��}{w{j��{���wv����3�+v�gۛ��3�����T��z����G+���2�F)}̉�m�= �nn�ff��;��O��������;�ܽ�v�=v��/�ˮx�5k��!���h�#�l�$�"������?��/�c`�t#K����]��g���v;p`�x|�MO�Y��iFEIڎ���A��p|i 2<���(�S�	JS��%���}��j����	�G�,d���o�6q��������z�*��@X�٥�=�ʕ1��j�A���Hު�Bb�����E�%����vw��l7�3?�3.����ܛ���%/y��:�L��$�i�����曾���,�p�n��[�v�z���v�}�:u���կy�}�3�q&4T����}�|;yO\���K.��Nߴ)l8q��s�MO��O�6O�7��2f����_��?8m��ɟv�<�iH�7�LyB��_�Wx`�?��?9�ă�҂TA��y�ۋPJ��߅Џ����n#;Ƭ�+[c�aL/<ݦ�o��Ҍg>̼Iq�����2�k-����ׯ_�M�G�ŵQ�g���?ӌ���_m5�S�T[�en�� ���'���ݠ�E[0'�F1�jں��v�E�:�Ǹ[,��-[�Q�
-e�(s]�`�5C,I	��N������&ug?F�׺g��/�T<+מ�C�=���vn����v�Y>�n�_��z�|�]��gYex��=w��w�9��[o?��;�ߖ�eY�� �w�9�������~sP�6�y�������q��yN�`�n���l���<����Co��%������~��=Ϸj��+H8���˗���rVϼ���#�i�U�]��:Y�x��+x7X��Wng���Ă��O���al�K��O����P����D�"����$#li�k=�T;Վ��׿��;��<���h�b.���7�5�ގiN��6��;�!Y��?����:��I����|�����{��p/��~�4�=��kҝ�|�@�����پ}{=�y�w���G\��ʗ�����}Ǩ?w׎3��;�<��;��?�C}� �E�۹ABŐK��G�c�6���[�G�]Dܻ���1�H��qr�?��+|s\p����o��B�F*öo�#�W��'�#��^|O���U2���}���X�QQgG�qQ����;X��X���y<��@L~�B���/��W���7n<� x#�g���t��RGS��ޜ�P�R��Ơ�S�Q�������)���U�:Ћ�NS���R�S��K�'_Fp�U�ߧe(�q=�+`KcS�ԗt܊9�8U4F��\i_���VAy	i���K���{�0�]1��$�-E�g�]o�]_���!M�R<���)�{����x�����FYG�N8�`���-Y��F��~���'7jYs��~ʮ��s����w<�~�g��fP����
��D֭Y�$�y��]�ن��lٲ&m�6_������7�j�-�����i���V�Pz�}c�\�R�tϯ���Ŀo�K0~��o��a��}��y��m[��������n;q!��������o��o��s�d���q�ڵ���N?ɿ��� -Tgڡ#���U2�p�dxdµ�4�9�L�D�Q�����PM�1���o�#��}���چ��tɪeL�)��C_S�_DB�S��X��mpe=��V��-ՙ[��{�oH@EXD��h]I�����ا�`s�*�w
��whR���+�9H�$���`9�+�\I�y�{�1��d��4��]j��zi�)Q!s Ƣ@4�W���[�S�I�и�GR�b�$��3�-%|-�豸�Z�1�l7ݦ�Y۰q��E���	`�;G��ƈ���6]�-����� �R���zd}���&����w�<��mXw�{��fBok.���M/�[ȕ�H�=w�m?��W{��*�Ɲ�w�b�y��v��N�d����XU�K�e�����AL�Ng)��г}�ͫ��!��0���P�|����M7�@�\��?�zB�c[t�l���=67�f��#G��<'���I7�E͉<�}�o�o~����ZǦ��m�HSɑ�BL(F�}�V{�������	�KlzpP��L*��L�k��"h�LQV��T�Y�.�g�E]��p�&���̝b,��k*ً���J��q�͈HZL��k|�Li&iD/M�O�h����x��� A�&02��5��B�T�Q��<VR/�TkH�N��1����7Xn� j@����h��5_Ms���'gё�Dl��}b�<R>SWg��᣶���m<:��5�Ǖ�
�7�%Y��esl,F��x�nإl#�?s����^�B�LL^9�8<S	���Ӏ�����`Lh8DB� p"dAspG'�"Li�R�r�'��e�(lT�c�ר7|qt�I��l��hZ,��TԴ�js�Te���{���[n����]WP���fQ�vO��g-��ZN����:��)T����(�ry��<L̉���� /$�|��y����H��d."N_qW}����Z�n��!���<� $�RB��M	�E8���ko*���I��N��4'��X�����ԝ&RK�r�W�%MC�!e
),���1�=�\��z�l�E�b�������� $'f��	��>����^�֐��]bip��A�RoTAEiiG�=e�;�:M�N~Xiv�V�]5�o���/�|�ݓR�M�W���B��ֽP{܏e���ZexT��4/���+?��#�#�c��9J���p~p�云�1��83�%�R#�Sw�6O1!M
B�u��9.��lxP��'��i�R�#�:b��G\Z����uu1HC�l�m$�[��Vk̅��݃�f�N�L ��}�s~ )��я~ԋt �����A��v�o*6�b��Z�0�9�	kRM)l�E�6O`R��3����,�v����Z���~�C�f!ց������)/�ą��`�}I׸Ѧi-B"����酂t����m��B4Io�1����N�s%�J*�4-b&��S%u����MꛘIJt�0oiM��_f�#�Ҷ`+����]�D�G�$~ER;�'�j 
*�I���<(��>�K学��Ms &�{5#����2�*�Ij[-��\��z\n�|��*�z�o3�?Vm���p���̡D���I�@/�������Jս�0���g��?�^���\;�0w����m:}K���@V����"i�7n8�?ɮ���c���K�4�{�C�	O����(�b�*�/�����a��g���a7���xҬ	� 'ok�֨�C�<b��[�T�3t�Dx��Xt<f��Q��~ac���\:TIWS��h��S��d±�y�c�
�]��6��Q�cY�T�f3��ii���`��}�K_r/ ��W��U����&�w�Pe����J�]�����T�?H��6R���C��ߒ��{H�ZYkŜ+�j�7ˈ*$�H嚛�r3����G�eҤz%��1N�2'1�h���~�.�`���UW]խ��/����uBJ�L�((�)�EED^k'����:i.S��bAz�$5�ߩ�Ͽy�~`��I���٠��-�l�t+�Dx��O�.E���ͯyJgR?��x�N;��	;p�q_?�w�w�%�������1�o}�[. ���o�׽�u��4^i���K/��|��#���5�"��g�T�u�6;�z�ӂ���iB�/��밖-ըV�Nx�?����k�,xp��]jc#�b�G��l�c�mzf���IĂ���Gm���v����!����&�j��w��~�w~� �R6��H[06� ))�F�֢�I�g�B;��KʡO������!��Q�����a�b�v���p����GV�č����
cÞ��s�׀�$127�Œ��\�P��Qaih|ǵ�G��Ԉ��#|]7���o�%�{!xz��J����E?d���r�|=�S�O�+���`v��u��������������g0~��7��>I���h(���d/�� �J|Ιgx�D���%H�h�A�i�,A]���>BK
ӉQ��@�觠4�*R�+���;�Rږ<���է�^�Do��p:��"G���O[����'�l8��k��f3��2�g��U�f\Pr�𑊯K�:���^W�o9�1����Z�?4 #����m����{�Vu�"��g:���6w���5�,�5���k��Bb'>��dtc"!ި��}�s,$��7o��[ny"0���P��DKk���?�.}Ƴl۶���1(P�߯l lr�5�4��<h���җ��Ŕ��2$��C��������=?d�F�8�p�5'���Ӟt�8�� �>�|�x"�M0n�'��D�&����F�ĀM�
��� �,�k9�h<HFƆ&�!๤��`2_�.���H��@8a��%!�-�l��!A���]|�Ů�+�"̞���w뭷v��@�!>0<�R�qE�h�It4�����A�!�`�3sG?��O/��wa8�^�>�����b#���@���x�'�42?ϔ��{��W�H柹�H�x L|Ƽ���\�#&s��A�b��ꓰ�ZJS�N�0w��&I?�S��A�EO��Ko�f���!.j�x��pK-��?g�N�jW\~i83hay�T�ߛ�eU2�ļ����3c2pb4�����e��A�0Rh�'���a��O��w��q�96_mط��M;x�q����Ex��v�%�k��,n�Z�;�;��^O�r<e^Nx�?����G������U��~����g_ye��Sv��ٶg�#{�ə�y��~#\x���áYX�S����1|��_����.���ȒhW6��5�yM�����Յ�-�����;ǼH�R!˴i��G�.�wo���^0�Xp:Q*,"� !�^�
c��"������5�saTC�s��0��I�A��������"9qX�~�p��< ��%X66`'y� ������Յhn�
qހ���?��3gR��ŕ��<�	.��ox�"am �H��ƚ2<��t\��[�������#���1?�@<��y6��y�X��w�ß�e�!в� �0�J+��z����H?���v���B�w�O�k�����ؙDj��Q�`r����=��nl0"����#�´��5�����9F�Zj�Z�	`�3`���;��EO;;G՘��J�8{��N��w�+~�5��.��מ�c&����?��.�ǚ�ߘOՕ�f�\��0`���c����]g�sٱ.���m:�p�+�a��kk�m�����H�n��˩
:��ۊg�N򖺖�0H]_���H
�2T�3w�gO��{�F٨�����t�MN(�"/!#��g>��@��90��]����)L��r�pl�E�ߴ�Pζ����*�@���ߎ�����+�(>$���VaqK��vߧ���o��*t�&O���
�8C��$^��A��;�⁔L�(BdyLAFK�ć�a <��z�R��?���l���BX����ε<��5��v��F��Y#�0DBȻ �Kpu8D���BZG��`\ya<���0��������\3��O�`2�����D��HPP�l*�Ë��H��^�җz?���Aq�����{�0�fO��y.�/���ó���jg^�/�m�� `�E����Fgh��"L��+���6�����Y�����A󥆯kP�6�`tl��ȯ7�\�/ʈ�%{��Tm�V�9?�N8t��Y�.�I^Br��������������~�;cK�N��g�3�v��}��b�]�%g���Z����O���1�+�aܴ�Ȑ=��>����j߻�6{ы^�O��G��9�g�a��c7�tC8��,I� ���w��UY�j��s?�sV��!�*�� ��QX�b�= A}��a�MR�uLK�(����V���A��s��˭��ѱ�OYA�ѹ�)o��֬�����F�5}R>s!� �8Iud����XUm�[Pb�D	�n��B�!��`y�C�3!�H�D'C����P"�qߣ���2�;#�N����!�2�)]8G:r���C��L߸��>�9�&3�0J�DzN��p�Xb���s��	�M�%�^�s�0�7�=�C������ɷ_�s�b�g<���	k�>��^<�x/ϓ��o�2��I�	�b�0��K��cXZA������vػ���;h�A�m Q�2b?���zw��w�c4�GZʾܰ!B{�G�7�}��Ky96�x��}�S��=�G^`�}�U~��:� ��e�Ұ�����/	�Ď19=h�Hē��q��A_��t0٬D����|SOL�q)��٨���Y��h2�	��|��ԧ>�Ź9���/����!X�WR�F[�7�����4f\M�b��P�e��@�[C/�\?Nl�O��6���B�|持��Ƈ�-�1C�������i�E�Q��q�H� �����ġ��sИ7��?�Y;�c�c.!�<�����!yq8a
4�H?�Fy'k!�O~+�C���x��$�2E`ƉF�{H�"��i�f �<�>\{��A���5h��E�1a'A��11�J���0*ր~ ��,	$"<�*#3sGc��H���a ����z a�AE0C��z�C�!�\#{�y&��z3_�����1�^�g���y�1��D�4��=���RD�S����΃�8;�By��]=��X7[� Ͻg?�*_'�L��g�9��=	�O�T���xff�v����n����Ӄ���Y��F�<��Y\�"��flx��t9�?��~߳�D󲯔��=;�+�y���^��9{$��#�_t�i%s�Ң
ד�&F9n���F�!��� �>�tH叾옺x}�vl??�3�67e<t�>�ߋ��ƭ�A>k�"����i-Vي��ϟ ,I���!��������!�G��F�c�:$Y5{��$�#�qCp�	`�=ćk!�ZS�!}�A�a�H��%D�y���_����� �a]Xs�v �:�4�OZ	?@9����!&̌�A�!�"���7Z��A�Ȣ%HC�9���� 0�����|���<m�Ly70�"M�^��k!��+���yd 8�Q%�A��}%+c��,����� ��|�o��~c,�V�j$�Ѱ�ܧ=���4�����4z/ۘe��y���u�].���gنM۬2<�I�b/#�gj��+:=2�| ��q��o��k{�A�!�1��)F�zMI��~�)�`����>�/0�=Q;�d���5������(�,Wm~n�\�s''��t�B��j1���/���
G��� wN��������Un_<��a�(�9_@9����u��D���kn��X��H2T��Ѣ�]�ɦ�v�7﹉���7<,�#�Qp���6z��J�Æ�@@88�D��o���Ɗ��R~��4\;-�.�7wfȔ߹����bǏ�R}����ɯ^��I��=H�rߤ��4�X;�ʡ�����s���> �L��&O��B�e`�/�[�ϣ�a�`��H��	s���p�>6�'����8`H�M��ɘ��O���y�x7��0�`5/�$�����\9�3Ew+e����@�����r>�qu��b���bzs~
���s�-�	����
�w=_�s�G;����ԟ
C��>���0/֗�����U��4'y��Cl�!ڂvkC�[���ͷ;�w;��ʼ�|v;���saP!X$r�,�c�Ĺ��&o�}���R	�$|�vb�W�h�4F�_��_�_��_w�3�� )�.�_wBɁH7��4���6:��B��!�p<���hƒ/e�7�"�|���4�q�����%��0u$�P!6V$b�{�l<gy���&�<宙F��^�S������C� ~��ȍPy��8$qy��7����lt��o���~����l<1�5�
L#�%	�@*��TiO��f>%,C"?�ٲ�X#��wA�h�B#A����G3�Y�xJK�z�4!}��ZZ�����$Qk�5W\�����8�vC[��J{��-�xK���.��ՊkQ.���z�������u2�	�ŹG�VW���cǝ�9C b_)c�������,h%��w�P���S'��-���\�K�nl��|;$�%�˝r����+��.^��|�qCG8�������A--�Ghg��)
Q��7�#p�x�B��</���p�W�Y�%Q��W��8D��`�N&DCɺn��B$0�}�E��d3(7��i~������o�I{�{�c��G����R�$u�ͽ��T���b�NAW���{�*`2��s�/��*	Sp^%�:�|�HV%HS����yz�,W;��
�V`��1�*xP�RF������� $��Rp}�s���� �Zl`�@�D��adozӛ���4��3�O����f��I{�A^\#�V�z¨�c:�2�k��'��	��0V���}���|ݫv5�5'�@����S��BA9�b�.@i�n3Ȝ�3cD�~P�.�!Q�����A]��ix
�ت7�}���2�6�n�DD*�?��So;	��V*��({����B�|'���R�ͥ�\њ5��� ����z�U8$�T�����ẇ�k���~w��˳GH���E6�.�K"�px�T�:b��W��'�nY�`�R�s���L۝�H�TAD��0p{��{�ԩ�5�D�%M��Hʥɏ;M�JҊh)���4�l*zF��&��RI�&��&`CW��O>��VD����oi�`�A��-f��c�g�)��h��]ஊt�D����ް��w�>1=��T�M��2"��U��[�-%���_o�~n��-�)�c[��3�/0�@�9����p����~��ֶ�y��M�f{�c6ng�n3˻&�7�F3��U���� cFg1O�W��񮶃���张̢0E��R��e��CY!�N���2�b!~��V��ϧ�+�\�&��Ri�Z�Z�v.&�r�' ���B&M�,Ҍ�:"N�p�5��:�{�����?l䃇��Ƀ67{ت�S���RD�$��v��5,�)d�I[K���?�%�J��Y`�TAT����q���H�H����C��xC�O�囘� �x�=���E�щܐ�	���&?�7ݣ흤�D��/4lt|��v��*hxl�S:S�	�A��k�-�BSFtN��i�i���\�f@�C����w��#��Q𿛭�f�t�
O�v�$5�jC�Q"m�W��w`�O�V��b��XʱPT*��E�)%y��3('�6-5�*�w9�Qj�l��8���x��c�Xo�@�|� �/dϴ���$��9��)#'������ϵ��q�?��=1�����sI������~���o��0��1�H�T���[;&v˵�-aM�%f�g�=�����5/�a�Uv�}�&�gl�m�7F���kڙF�g�`K5i3�UE���������vF��Eo�J	���\����^�|�[�J���d� $��m��A����S�q@�C�OE�e����� -2��S�JM�y��;���}���{S�}+��V��sso��9�����k���n�bwio�ji�I߽�_�w{��٢!(�8� ���=�y�8�Ѳiy6A�u~�l1���g������ ���o�׎?ꖂ@�y��`o��2"�ԭ�x.\y�%>c�����,b�CS�y���t(�"xMj!�C���� ��$E��ԷS���(9�QMk4�b��?�JX(��F�.��U�U�<���^z1w�d7�HǆJq�w2H�c%k4���)�.#F���2{_5�q�8/�Kl��٠�F�c.�[�,�1�[��[¿���{r��{��l��7��1�胱��-���/|ZU�jH(*-3m�F��m.mBY|��ִ�����1���w���ش���5t2W�mgƎ>�@�1����x9W��C���p�F(���K=�۟�7��(J���=J�
�5��}�m����(�!C���H��t�8��B�^o��C�l�S'-�rm��6��=�l߁63�g:�X��ke���BZMk���a�-�6�e�f .5�[/W0���؍��>�Ϊ�1KY\����l��_w��h�:��V ��*^� �8b���.*}�LF
��C0��'UX�s�=ç9㔰P:C�i6\�ѩ�C���J���{�z7kh��K�t�ދGB��&�W �e#^�R)2��Gy�i@��c����<��o?RlyY)=�S)������x��V��xtσ֜���Y��#�{�68�4
��c�`��h��9�i4�jQ�ˣO��c���֑bX� L�3zx�B.�(���p]O��f�GP�L���)�8��ӛ���pH�Y J�І���u��q�6z����\8��H���=���<?o�*�k���$ɷF�:ַ��M�ۻ�����gN�sAX�mf�4�jA1�4(1}l��u��l���^<i�A�GDe��l�m��Yrɹ��+��t�b���S��!�I+!AB_�~���X�ݳx84ۊEu#�a�U�ޖ��.x4b��ʵv�78�?¿X�� \�ctXO]�fpl�Zq����e@�H?�W�ݣC�v����ڵ��l	�DؿȔ}���:~���QF��l)�xQf�g���w�7;�9�(���[��thb����@��P/FF�o�s���դ)r��W�RC�9�R`J�y�K�q���_�u�Ycf2X'eg�t�C�+�q߾�v��;���	+v+1w8�~�3T0Js�(FEX�mW�
������� T{0;?��� d�H��9)��;;��-�'Y�m��Mv�5��=��a�y�aC�5�޼�;�o�s]O�hw��ʷ��O��Wz-P�����W��I��~R�N�_��_w&�^�9�?ˮ��*۲ꐚW ǽ�p���;wy<�{��.���ډ3�+v���x<��z�>e��,�x���꫟f/�����#�7�b��N?A�5:u�t�F��M�(`-$ �!%�L 	w^G�� �����5���^¿ ^9i���A.�?iǚs*!�m,�ȩ��SA���S�D ���}���g
R������?�`8C�sJ�¡��-���6�*�v-�5�d�<=���`��V�����1���E?�9�I�����2kU8_��ʏ����W��X%��9n�	�Xj��߲ҕ���	�ѽWE�O1(UO�ޫHOך>�����T��Y=c���2�^�:lB/�b9X�e
9�� h�M�c�a�XS�x�b"����V���&$=��/���e=c����y���ʯ��i�c��q{�w�]�4z.�����0�i/Ɯ����aՒ]v�v�,�`�o�����OkI�EO�%�Y/��/K��i5���`�o��K^�"p"�v{����o���M���~����.��R[�f�5�mgy�RH�*Q� �P<7}�o�[�3h���^+�����"^�q�	�L}&,Jf�y��۴����=웶������8
����t���Z6"H�� ��Vo�TA�f�k�8m�"�Q	c�$�T���u�W�Jx��ƙ/sRe�)ǉy�Ŝo�!���L\Li1��sD�s�񚠕4Q@<>\�^^�x~�)#Jկ���� .C�E��1�7�4����ž��(w��n�����7��Iqn4fmr�v�jC��-Y
mv;�,ve�k�f�s�&����f�n�F�4�������3�8�c�%;�԰��:���S'�ѕg
/���p���k�pf ք�si"��9j�zw(w�;lF�ú5k�&��z���Лv����W�h���u;~���DXl�w�];�ˮ�:�k79.�u�۱#G�?!�b�r
7^���|�+_��n}�m�h�������Nu,���!�=��]�a������lf�D�\:��6���OeHx���={���g��>�����݅�;�����pg���V���n�
ȕ�W�]��x*P�P`��<��g>�Y'�b�_��BO5U{C�!�̙�1�&('x:<g�X�����wZaxpD�FM�g��5r\|膁渖ok����"(�����4u1?Xo�������q쑱Q_�:?���D��A��uk�z�0�����gW@w���p�T�)�߅bֱ������ׂY�z�:[�bC�#I���Q	�:��kϟCDn��0��a�Řbm.J+�e�8��m���{���ҿ��;��!U�q�5��u7��T3�^z�S~�C��1�J)M 9��_잣�O/˟��Y*XU͸�ᡟ�:IbU�����^5j�.X�<:�z���C��׾����v���C��!��WJ��>��hr�0<(�U~�'^�^	���C_�<X)�ël��~��{�}v8,".��N�F���cq�g��i� Z�<6@���kEB��B�@���?��@3 m3��=z�K^����@�c5!�9��P(T,u���a� ��)�a�y9���պPMVd53W�)�!_�� �Ie�o���qm(+<<8͕ J��v���p��;�A^m���C`p?FǆGFI��������X�Pf����7����\8�ڱm�Si0w�k��͚R��<�_o)*��d�cࣣ+m3m��(�f���n,�,,��0$`�Ϭ���W�Q$cH-�'���>�g�� 2����e�U�ׯ%<�o�sή��
��w%�F���O}�� .��i��o{5��?���v���7����/�3X�q��:��YK��_����Um�u�o�� �&�R�88¦:v�MN�� k��M.��x����8�#*`�QYs����y
Xt�z)��u����EpO���-�u� XA?p��V0���52~���;|�#��H�r���2E��X�m'����~�y�#>���ѹO|���� ����[�l��,�Ga �x&��s%���h��q�5kW9$ǳ�y�]~�����\�q|^Ûcsc��9#����(����!���k�E����-QT\J��̱yM� mjR�|)�n��5ǽC�n���Y?NW�.��Șٱj��{	�V����q7��m��I�J��P ���{�)T9P��s^�a�7rl�F
=��]�z��q�����=��ɣ��r1��k�s�3M/���b�䄑X���������.��a��+��w�;�����/���gݶekx�-k�j�#��7^ikVӏv�ff��=�`eWmo��4� �og��+M==y�~���E�B~N�K��K�sW��)q�b.�^����j�����>�KG<b1/}��Kv1�VӨ)����'%KU�(�#�Dt&FL�����-�"����/ӿ��Ω"�p���J�yFT�JC4'������;Ne2BQ�Xxfs��~L�;׆���t���N�^���nܜ�&�0�3�=2=x�(
Un�lX�^tA @����}�QkD�+�{3J�/�>;���ZA` ,/<��銻}��6;q�S�[(D"8h���aO��ۥ#v�nŘ�O])��)���;��k�u�4g�A�¡ D��*>�z���Ԥ=��=�rŰ������#���v�G�R*ة'��ذ�B��}op^���z�g� �z�_��Rtv���XN��� �N�,����a�@fV�F.�"��v=h�a���dP#���Q�?��?�M�Pb! U ���Xo��|_��d!(K�x�Ҋ�Ƭ�*0�6�њ���ɰ ໯�p�.gt+,��l�B�yh������]X� e��������X�,�f�����P�\;K� �5&x*J�󲱸'p�K�=���~,0��g~�g\� ��g��fR������[�ͥ�s��=�v��
�d�_6=�k��g�ry���kF�?���v%����'̕��@�̵���kc.bC�U3z��2a]�X�W�s�p>�g��1pϸ/jCyn�QH	tm1�?)�<�X�_u�W ��=yb�V��|��6�L��I�pK=���l,�6/eee1�Y�@|�4s����«{��{l��Ƿ:�g�E�p����S���0�B,���W�<��̉���?�y��IY���(��̔oڑQ6����A*�U,Kl�)��iz�f#�T�u
f~����R��y�b{!��c���9;tp���}oX��66^��k���E��@YZX�۷�#C����+A܁�@F��E���k\/��DM̱���5���N"�k������:΋@�;Vp6��c']�#�Ԝ��،��^����.3s^�zE313�XPףt\^G�)~�@�o�r繂���|��Ԁ럘��������Vf���G�P&x��ȍ�qn�w��^
־�1��	؇�T�8��i�FA�5.͖w�b�;~Ć�ﱡ�UaM�[��{��k�#���S�����
��������a�������7����z`Ȩ��Ӛ���ke�(z�d��"��"�@��b,qxd��Z�"W,O�"���)��>7��l�]]Z'���Ց�)~=��K�r��[��7l��%�V��p[�l\�����?�������\y>wki^���e�?l�sAIET�3g	��E�(�"��ur�[͠h,X����u�0����H�s���j�
V��/pKA�2�
e���~b#x�pB8��`��^�ʯ�?~��杺���[�¬1W�k���.�q������#�jժ�֨ovܡAM�/Ͻ�9. 9��ب7�n4��ޭϸ�ߓ"`�dg���}��ܺ���+"$�7�.Jx��5���O~}ܓ���%�l|�F�m����k,���~�w�r|��Wlz�7���;��B���r�����(��[�9d�<Pd���/�y=�Y�v����� EI\��0/�~AJ[M���<U��0�RC��& Ȱ�qTӡX�֧��i���TťF�!���� �뾐d�p�[����xk{k�T�e��1[��v\r��׃< #���S1hɕ��q�Q�����[�?��'��\د����ۯ�����ҋ/� �����)��JT�%�@���Q�t#�X��t-�W�@3�ylx$�g�T�K���R�y���j�W�!K;���vX��9�k�{�iG�����w�k��9�U5�E����ի^�P�0ؼd!�����j+&�Q!m^64�D���>;z����e�*��$T�˖�B����Y�g(�
�m{��^
 �}bO���0	N ��և4����pN��9�Q�/֋Z�?�wP��,&yBx�2�a�s��fD�'�+X��u|�s����C9��zZ���1����J�L�5悧!aԣ4���f~��c)5��B������.�E2o5@W<F���Ҋ�MxWR�D�K��X��� ,]JR���v��z���PŸ���R�.='N�f@�3�^��sL\����(���8y�{�T��'�Z�S��k�(_������B��~Ϟ=�'�'��׼�[���-o�,Ω&���W=ﱆQԫ׭��bSӳN�7^̮ەV���ȕ�e���Q8ݵ�Ϡ�Wp��b�7��W<88����_���pݵޡ�۞���C�e0n���uހ�߰2<Ԫ�;p̨�A����K��y���wz0\�\v�BXW]s�o~`m�٬� kyfz������f��m��a;9=���iD��r\� y�r!�+�y��~C}dU��o>?���`�"�����`��]�U5C�H�_�zsU>#��&���yO�T`�X��6���P�����>|�M�5�y��F癨Z�g�޳�_躽7l�M�1���|�P��96�������ؐȫ�[V����^�PR�Zi�8	"Yв��B�@SN��	�*ӊg�ȩ��e��U�:w���ɭ~>j�����c����W�Y�4΁�H�H%& v
���DY�z���H�W�4��eu7s��\�X뭬��@'�?��'&��|���.�](؀��2��=i�&gmhxܠsvt!�Y���7���}�+�؁�/��灂�"Y\��H���"�L�.9�Ë}߽��ϼ���Y�x�6����AV��]87���[��E���s��n8>�?b�T{F�Ӽ��O+6�!��bx������+e�ґ�>�屑!۾m��_����:x�<�a����CA��=�U���BV�������.�!m��K/w�W����&vh&\#�3B�F�@{�	��`8/�
�C	�0�xE;Q����3�u)F�2�\�36PP0�	e�<H��~��x<���o|�=���Z�(pu��N �{� g(�����q��|�����/��9��F�=�<o�d�[�� 歴����=���=�뮻|=)�V7K�˛J!��}Rn����LxJI�8��RPEw
󤰍��������+�,a��+���-��!�+� �=X{����_�����a��iZ,�g�'�{�}�^����~�����R%�ͺ-�o���@x���<P��Y�����u�:�sb �Y�x��o��M�k��|l�~�k����4�A�tl�m�y�%���M604hS�s����B����g��_  �f��j���ȋ�O|���[���m�~�w�yd�^۵�A����+H���˞f�_y�]|�����qc�k��h��_�W��y�L��E/z���%
�C8h#�z�ڂ�ynz�>��OZs��!-��1����5@�<������`��]R��+��źP���z�k_���?����� <�������T4 
�J�K"P�%������Cyb�*�&�0L���tL�/�D����gȖa�!Xو(���o��m����i��{,8Rq�\?��?�0X.�h2}ڲ�Q"�x���.8���T�F�=YK(���7��9���7�1���^ )��e��%lH��f@�Eֵ�q�P��iuu<y6�w�
l�C�N���dm��.VZg2���{ �y-���?6e*���ݳ��{����A91��-/_�6+mbr�ceP����;mF�����'�vvO)Q�C��d�Gq���+5`X7�x}�C�֭�b���>��]-W|Τ��_�=�����z�&��a����g��q�q��~�
ݚ o?˹F�>��Ϻ۲��`��ƛnJ�{��~��`�+׬���.�e�"��E� ���ᘈ�������rx��a��Y�A!�$��<��wx�w�=_����`��:�!�(�u>zl6���rh!�Se/n��>�-/�1/��Qn=�M��MДkG���6���Kγ 12�E�	�b3pl�G�V$���*����̅{I�%n/
��3��=�H���B/�����;��fnT�FOf��/ރ�Ұ�����`����VQYH̓�^k�B����O��	b�S��Ҩ�F��'� ������[ǂ�u,>�='�h�S���1�*W	qF��W,@�[�B0����Q�<C�-o�����[���ӟc��1[�r؊����ʞ�I�;�=�5�6���yn��K�o�} yld��R*�'�w�?\�!��M�X^ׅ����FQ�$���Xx��֯�U�/��n��[w��?u��2��o��6m���0�w���ѻ?����+�Y/��ֻ�;�T1p��`�~d��ٟ��^��Av���k�k���HŬ�:��X�ln�VA$
�)��`RV�\������tK�E��������w(
B����Y�Oz��T�f.;,�/��S�V_�e1  ��IDAT�9�N[ذ�������
��=��3�&�
��,|\�T����@�\#�8��1Ҥl�(�
!���Ȇ�ް�8BOE���Gys��e�f�R�����h�3�g��E�rI1rY�\�,e:�����~l��!�Y#|��B��s=��ǣ��Ul�$DdK(J Kp��K(+� ����
�+���4{DB\i��e����|����$#�y�K橸�2�4o�)-EvU���n�Ev��WS�y��V���gf���[��+lj���1�|h�X��O*���tO=#�򛜎�is�>g�췗������~��z�Z^EVpr�{�����^��^�5<�<X�+l�E�mnfֳ�FG��.�+~�#=�ȁJ����9w�8v{��O����N�� C@��Y��@,�w������n��6�,V�ɐi�,��Y��>v�G\`i��0��@����q���Y��=�x�;��X��%J�%1#E5(�JǙ;K���
E�}
��_��]gb�D��oȃA�2#�	sF���#\�����pl�9� �V�ŀ�&�{bGDx��;���?`"e�7/�����: ��6B�\z} JE�[�����r~�q)���
��X��^��;�c.̕�t���qߠd�C�,��3PSp���|��ZB9W�U�Pe�p-|�����P�fjy���R8U��"0�#�B� ��#��*��uy|(��� ���y���k�xf\� ��?�A���c����8Ć���}�T����U�"��{h�f�Vۋ�ʵj�������E��@V�u(F���5�������]D�X�y�S�[����g]��-��]���62dM0̠�����=�v��G?l����3�ckiI����6��ހ0�&�ed�<�QK����}&XjP ಣP�G�G�Gz8,��f'���k�"E� ��q6�d� (X<��ۿ���i^�R4�u]YMMUm��	+���κ���wߧ��r�c}���c�C�{���@8^x�_��}�V�QH�D��9�"�6 �S6,��������TF�
������
G�1�!����B �>�dc"�`׽��r.�P%�|�7�e����>��7��
�p�@ �!�U�P�?�˵s������b`�PM0W��'k=%����d�=��FW�X�y��,U/�kn��V��ز ���Ǽ喙0�geYO���{)���=��e8ʑs��Pp
��.�4뽖Ѧ��R������_p��l����ɪ����2͍���)��[#��s��ǗŶ�@��Ś�B�}S0&/��J�X�������͠+ŮD�r��q�����,�L7���k����` pe�{�.?PQ�9�5 ^Љ�]j���
��?�!�{��͌�˩�x��	�]�ͷ4,��dq��45�ZeC�`�������/����O��
,�3�����Mn�⡽�>,�^�V+�>��.w���-.��5d5���E�@pE���:x�+_��닻�)k��]@����`T������T����l~��jV̣��:J���	kW�+c�%��W��7�r�����ͼ��:O5D�U�&�e{`щ���'�'�G��֑��T�(�+����\���&����J�w�f�Q���hrr�_S�XP�j�Ny�"!�'�|��"x]�(3k���W�*2���L��u�
��B��_R؉������kG	����5����J��u�&[�vC�C���F�f��2Z�ڡ����=�p�IH�0եp�����T�Ǌ��=���S�>�;*ume�Vx
"����no̿�]�'�]�5�e��Q24�7>ZT��B:5�� �X>���M�<��M�Wit���k��`�u�b�F�����Nc�n����pz:����H�Q�
T
���B~��2L�`����� ,��?P,@-Ef�Nf�7i����g�0r�<�ShcJ��hKA;s�ֲ�����"!��+y��z������*|�^H8����dR�^�J�F���q}�#c�-%����*^W� �3�,87�e��=��o{�E2�����`�c�
�K��p������\熍�eW\�ﱽ��t���=�����u�����f)�<�/$,��"�U��i��vs>�薧}�+
�#�?I���_z�Vw�����g�#>\��Aq�U��ǟW�]�٨��+k�_?���Ŝ��=�=8������xj���6gJ�Y/����q�t�eeҼ��n{�MۚO�K����nXWX���z˒����K�Y
��z&+����)g�B��Uv`��� )�>�8�AX0X&���gr\�,P M�N,<�U���lp,HÁ8��9��8J`#ă/���p��b�*$��=T�
�HlŋUJ��x��z���,�� ��9�I<�(���x�9�+׎@d���/!�g�G���cP2 �Rذ�|�����ٟn���z3��7� W�UB!�V��WU��2uXlz�9�Ph����
v#��\|����s.����꠆ף �<�����j�9ǥ�u%��5_���+��ݏů�n�#��9�ei�Sa�<��=�z�Iߠ{h4;q��b@5镲 ��t���)���?�'�5�<P*ts�گ��BLKu�"�X��sc������_�a�g�-�j>�E̕@K$K����<�����))��=<,R9��~�^���yF�K��#�û�M-gF�5�"��W���^2��,�Y�W�&��{�U׸ %�K�
��I�;���{�\���Gq�7	���0J�+��Pmx����;��L}�
����h��LP4�B���rl�N)�B��CJ�� ��9�
����5��X�j�5�f�w������,���

�`�ū̚�j5� ����x���� +J���2�!��0�W������7����1�N!�̑�@�F�P�iL(BYJ�-o.b�B�F%��'���y�*�z�b&��B���S
�̯����ql���(ԭ�l)�<���B���VF���4+�LZh���U���`�n�/�p��m��gPP����c�I9) �,��^@�s�e�� �2x�E�����F����������p.\�au<_�=���l�ѱ�3x�:E6E�S������M�/]kl�"��d��ĺEp��!���۵k����w |�4W�늴J,o�K�t	*	8��c����y+�4B����_A��H�D��u��7��F�� w�X�j��2R�s�-�5s�(3���ÛA90v*��!�D_�y�����+~e�(@�5�I��$P|�&�7����hE�Y*�|xA�?���\��E��d��� �h�����Y����\}��2���,.%υg�ץ���'��f��ĜQ�<_M
�i��"�no/6�]=����Bs�p�C��U[�:�̍���9O���Պ�n�� �<G}L����5������T�d���h:��E���0�b�9Z���?�������9��3Y8< ϭ.ƻ�ng<&����Sˀ�|`2D�'#b3w��  �c�%�=�J�;q���}Ȏ���
V!V6OS��-�O'��S�TQ*X �4�a����Z�H�!@����4]EFlz�� .}>�1�TʒM�<��s?e2�F�qQ8X�X� U_^��\�x�;�ax��L
#�J-�\��5�=�X�y`=��B��� �a>QAY�YLɬ vz�h�z�:Jc�+u%���c�O��&��5 'I!��<A�xR�>���m�>�_1Y�xO�o�פ�Vz��I�H��!�J=���N^���w~�b�b[�Jl{X�1��	*����.�r�_#�V#��Y+-��n�'U���Ih����x@�qnJՍ��R��]�օ�g":����3�.�g���������6`NY�-��}ou������W�7��).o_�5�$ L���m��p
k����c�lr☍��j�#�2�}��+͔�gyZ�!��<�����o�'m���%s�_�`�>��Kإ�����"l��:�G>x@-�!�!�KU���e��"�
���!��+���%��2��`05������ �X����=�n]*fJy��kd�xR^�zRПav����L��!��)K���K��Q��k(t�T����������ͣ�"�w���3n�նl�(�����~�a]�ךd.ɂ-'�l)*��g��]����������9���٨ (ҀX�N��)���nVx�S;Ik�">ǉ��{[��	߲��4��h�W$ռ�Q�h�~�w�x�2:a^�v�;�6�E��_7�s�ȫ7��r2��S4[u��|�U�q����NA�,�>���i��$�ѣlwb�03�T��5����A,���p^]y�l"��XlY}���V�v��c��J){Eo!,�f�b���=��٘�e���@�|A#�a�#���������6� �p=�{ѵ�]V
!&]τ�c}�#OP% FL= ��e ����Е)�Fձh��|�ǀ@�~S? U��ൠ����|AF���I� �@m�><M���L�Ac��&hG�>ץ�]�,�@x��s��f�(0�BF��f)\���0�fI	��N��Z�����ܴ�����~�ɩS.\f��5W*�zZ\�
p]k��n��sn���W��� H=)6�Ou�4%��$:����t�3���m;?W̕+�
��O���^~���-W�P%�ً��'B
u����=/�?35�ߋf���������-��{����F*��-pE�9wP&���t�)���9�X���x}��۹<
���k9�D������4#L.ndi�ܞ�8�F�"��z-���*���)>����^B?��+=u=a=zd"X�E��� h�5�A67\�z��Y(s��7�6�(��SgScR��,0	8��.X��M������0{捀U����P�g�����d���je� ���̊���s`�@7���~���>�<��96��<,w	@��T�)m����A�)�ϛ���R�����86�'�+�WZ�80��ԪR9�R�R��$,w\�.*�ytM�:��w���o�-�̇�������yC�c)���3�"D�\�=�}��
�����kIXCs����y�
r�6@���	�[z�L��,jf6x/��%��9/جt�г٘�}�w�Z����>׾��1sϫ���(dJv�R��f����7F�e�s��'O�c���#p���-,h��N	�c��Z�:�?����oΝ��;W����nӘ��3\���2F�%�.h��\�^5k�*?l�Us>t����e' א�'�[A1Ǣ�D��t�?�͖��x��a�
�xF�\*����U6[��M����d����[x��s��s!��p�4��5��'Rl�G*]/~�	�� �W.�R�<�e�I��}��bl�����	���X��A�my���,�f��EX����+�y�0�����S�B�_P����B']_��jϿ����#s/4[+��S�H�&��p&q��<#�%�;�����{�>	x���(���Δ���bAZ��պ��y;�W�$u��IኧI�N�������&[����{eͶ���q���M���N�\��{-(�L�1�b�i�펧���?<<j/{ɋ=A ��b^�������9J��^�g+�@c@"W)Ÿ��̔{Jp�7W� �9o�ĺ���q��Ɏ�_��������j�@�}����y�V�:d�@�w���BD
,|Y<
���O�X�T����,#B�-�������Q;z���;�E,�V3α)�FƖ�l�aC���A��#�U��֏Z��+g�4�X�??�@6�|^�b?�-A.�T�\�Y��LBL�.���\��#!�znj|�"2e�nR�+��\%����ϊHB_�A�H��o	���ы����(��*�!~bg�Nn�ׯ3:����J��/IC�&	e�-`.>����{)/����o�)����Z�B�����C«�d6q^���`z&�D�.�
G�NJM�a^��V�z�s���a��lnf�s����䐞��[6�Үw>���g�
8Oɔ��o�s��L��=�g؋^�b{�[���.�w���5���ZԞQЛ�B�əY?���k���$��Q��r�a�}�p��Y�7�Yz���P��*@���ew�U�r�j�`�\*n��_�����S�G��6��Y��cA�o	Yy(8����`�B�~�{�ч�e0����Y�B��g��{��y�a���K���w=#������x��k .Y^�Aۮs�p�'ON���H�јuET(�l�ju �{�s�*�X���l����`���BX,�
�!��Ț!HŻ�e0J����}�;((6��Ș����ȣG�g��M��S��>�h���e������ �v>����j�=�� �)z�(ޗ!�w9���k���0T`W0�`��������e M��DU8���9��;#��s��/���ۻ�ֆ�T��D�c�i�P�C��p��GF�TfAn����3J���V��@,�����n���Ea���Zv�����M�=�r������}ͮw�r��(��|o�˷9��1Q�P�P�� /�����(C��L�FO(���O:/��7���8
��# �Y�G���|���E1{	:���3��H�8G{�v�0$(����Lx#t�կr��a�V9��Lh�Ć��sa��'�&lU֭�>YK��L)�rs, �@�.)�i�2��j����@�.��V�;l��I���]1��`�ݒ�x��>+@�L���K.��5(���ov�"�2H�)��9�k+%S|/d�|�w=��X7��ʓ�(�����$%��$0xj��UK��%?�E�%@�(YJl.��$��&'<o�2!���,|^�:���%e �;�Y�E��?�"��^�qI]�>�*��<H�Խ��|��� �h,t�di�����}�(��	]�&�&����1��{��E�0_�����U����K+Wr1���mr_�kN3�� �'*ϰV�\�$�/������^h��2������9gqu�C���(���LLĊhkG�\����K�-˖۝/{�C��aR��c]��e[�f��ر�>����������A�]��ȓg���7�ǣ�x��٫^���za�fc�EK~ �~tt�Ɨ��-�0�*h)��1ɒa����E"�EJ0T<X�l`�}ua�9=.���W�,�bݩ��S,�4����\}*K�+�5C;�6��aS�ؘ󕅧�m��s��J[��2�2��AKZ%�A��M�~�(ā��E`Rp%:,Yb(A,"�K�'J!M@�cq.�T�у���TL�� �Q�(-�[j.�0`ŒWz(���Qr=	�r�Xn;�����,f��=�؍�B1�bD0���W�<�j�@��z�����
e�\"�	�4՘!�ε��P�j�.��X�֋��GZ4���j�Y����/��/�ڱ����x���;�d��������f��1���Pg��;'�,�P
JmOi6��4��i�}�I�+*��h�N۝�M5:��S�s}���� 2SN�Y�O�Ӏ��oϞ��>f�)���W����ړ�K�-�hX�ϸ�&�pi�hjjjL*/,c��j��9�U�8���)oϪ��Of���!�E�f�*�>Y�j�����{Ͻ���v�����Y	s%<��o����&o�c�E�1�"����&��g�gsܛ�A
".$.6��Rz�F��U���r��E]O#]�|u��5fO:��C>�*yJ�Sp׶P�Խ��W!��(�兒�|���UW�k���9#�j,N&V1����w�6%��M"J�h=E�%��EѢ8�.
��x��PЏ���pN	p6$B%�����h��$� ��s�������>���{'��MLsn��(R>U��w�f��1�dF�b�z?�M��:@��ޑ�z���2\R�����Q TEE��S�Y���KR�1��3KV�iv�Y�C�K��7J�NuY�:��KMg0�����H�����'ҘA�{�&&�����%S��$��
{�ہ�o���.'W�+|��J���
t�{�A��zXC����x���opo�����"��P��g�S�K���v��kS����#�/���o�kxN9Lz�u�������{1zX���G2���n��}��;ۇ����A�_v��v��O3x�[A�۳���_m��a۸�r�T���%���gϼ�v��W��@`�R8��J��(��Y lr�����l����-�4�s��-($kl��m�z�f��>n���¼���:O��w=��sY������a(���a�b�"���" �0X�@���{jW�k�@�3 -�{�E� ĺ>�7�e���`�J�?c�ca�T�~���Y���&eǨ��������� #��|�NA+\�j�9�h�sǺOy]t�P�<s ��84\B^V"
����?��� ���	�WN����ZZ���k�Z�>(k��9?���Ȩ��f1��S�ǳz��_�`���ՙN1
]�e/��4;Ią�����1�`���}���U[j��>Z���(���6ۚ���_a����C#nu:��V�I�����E��� ��w|��W�Ws
�=q��N[�ض��v�׾���
�t]�+"�i�БÏ����{�9w|��_����M7�b��~�ב`�T������/�����ٺ����M=����o�@�����8h�.wpjj�N��6�χ>�A�x�� A��sYQ�Q����	k���X�i%c�٢�z���b� ��Ҵ�e�e�k�7��2�x��0��sb���u��ӿ���֪Rf����Y����9?�!�U�L,{�9���_��s�4V5�� �ʔ��ō%����gs!D(�����a�X��<���]'X����y!��c�i����!��(&��uE�9�r�y�¶96�F��>����R��+HY7�(�aH�������7bJ��!�eaQ2�0Pe�}�e��:���a�k6����&\��;����2���dw���\�,y"��bAٙ�Ӫ�Փ^
���\;�|ݰ��s-��+�A��|{��[-��kT�chx�"kUƑ�Rd݋J�xz~$LM�8a�����o���p)��:�@��������W�x�����pҳ�%���i�w#�Y����T��˯��Ղ=���v�U��E�օM��Iϝ7?��u}:��e;����?�^���������\$d��ԉ��#�x�q�Aq�����¢��y�>z$w����}��[KV*EXyzZ1rxƍ���Ѕ3������rJGeQSEK�
x��d�ј�t��",��jD@#0�,BP]�Ԏ+�{�o6B��`�# �Q	�b)��S?�S���"WC!a�� Q��&���?ޘ�����X|�g̃2�k!��5���� ���>q� "`%�2c�\�ϱ��|��5A#d�p���)��Y��SS��+�eq�1�Tx:�JMv7/��%��En��o��1x�z�|�9I!�90g>#8�g�{|�S��g\����B���9e�Ⱥ��`<��G!YۋX=S�G���Z�زѱX���oY�V��`q#�wQ�ԝa���>��v������*������/��/�JC�!�x�x��`կ�fk¦�&���.yOP���<�^��o���*a��\����zљX���^����?4<�س;�s��:d�`={�CC1`Y���Z)z��MDe=��c�n8�?�s?�.?��B���~��XlJӫs:�?��n����O�KZ�d����U31y���3J�
�T%��$��9"�����H&����c(e���0 ���AEW|Ndp|����P 
�i��5`�r<��#�M-�2��=W�.�����w�����( )60J���#^�Uv�@H�(M�8�l�(�h="�Sȱz�S�[�4z�tXk�����=I�r/�)�9�p�0#J� �o��o��������yQ<�Ng��k����_��1GY�o{����\?�Hyf��{�r�5xq�K0���<	�`�s���y�y�]�(1=9�$
��cC�A@�O�G�@Φ�A9�xm@ ����܌�{NOO���
+Vm��q�dDF1#O�n+#v�gdU�&����1o���|��Wݐ�6�}�q�;d{v�
��B��jՠ���(�:k����{����r�3=^�^�:�}�b8Od����zc�1�]8��kqC� ��ix�O'X+v<ȄU_�2UySS'�����0p<��(����TH� p�����1�(-.�⧥�5�_D@O���ܢ'C���R�Y<cˣjV�> �P�i��;q���o橬���4�F�^}��2E8���%�l�3���6m�����íJQ-fq��`�����)}!��CmJa����b��+���ڎg�}q�W��ann&ǳ!��ξ[�J�;,L�x����q�V$�	]�=�ɿ�ï���9��������y�A���=�;�U�R�+k5-��9���y"��b�f�i�0w<�>���|�Z��
k��Z�
n�[����0��۰�yF#c'�@��ŋ뱩{��J 7�2���pY���`y _w�e����ed)u��g4X��@�4O�si��SB��g��r���}7<����~-v��n��
�X�[���!k7c~8<�Q`�S6��i�k�"��[��X�0KY�(�#p:0oa����h�BL@D��|���\�N��"���`���	�F��h6�R��4��[:��7�*V��)+9�#��kVPQx����̊"A
D�CA��V�Q�@�nZѫ�p\�V�'������[]��-*�Z̬�
`���ôЌ����֐�"�b)l^�󋋲Ty�Z~�P�������R�(�9?����MF��5�y��&���-�����P�����Z�x)�/J઒5-@C��$kIy���=�	����ow8�,1�jyF2���b(Z��w�M�ܵ���}�㠪�j�Ra��,8�?���G�v�X��Gl��N��iv3�:ˈ��N砤����l6x.@�p�?Yh��T��5�����+�jPp혵�=�v�Ѻ��1�Í��P��r�Ki�)�G/��y��!��y���d����A���j<�bL�D�V��)
5���c�P�	$�xpP
��	:;�!qq	b��>��M�⽲p�������c;�՜
�aN���i`�x;�zv���]xͲ&�=�(�S��`u;'��~	�Џ,e�H��yT ���:�\|5�Q��
�Dɠ@eJ��V�J���_/�%��*���)%�YB[��g�yu:?�PE����=�L�e��6���C�{!������ҌyaĚ�b�I����Q�T=�Y�7��ҕE�̓��	?��c����x�<��=R��A��ʘ�:ԁ}����K���"����}V��<�F�!�9� ��e��8Vu����X��O���m�v�� �n��w�\�Gcü���±�v���/5�W}�x��5���� ���(v+�2��ky�������v�8����������)���[zo�¿'m�,@��b��kæ>f�\|�ՃU276aa�jU�
�j��D����h�pW5��R�X,l򾱪�_���zVi�X��nq��M!���`��)=�}��F9�@m�f&OXi .��/D��Sh��螮�E��@#���|QG�k�*S�*�,��զ�q*�9����ɛ,e��m��;�D������"v���)��M+��{A*���'˞���NQ�oR����b���GE��x_�E�:X/BP�|GN�R'SG�S�'�R�j1NDy��!6J֯��xMp�FZI���EV����hR7�Eʇ���}5�)��ސ��Q
�7<%��p]��ĝ�_ۧ[���Y��X��	����7u��k)V���O>Go\�)�궜W+�Y���;_~��Q�"xU2��A�P��z����X�p�I�8yȦf��h<{otl�O�ѵ�[���=��9���h ���@����R���/��pn�G�n���%��+�28d;.}��~t��{�q�/�ff	tl,l�Ma��p�[�v�?��Nz[F���f�0�ʀß�?15i>������ٙ\�a�PQ.4��m"��o|�]WT�2�,�Y�p.Ulr�aA&��ȐMM#`��מ�b�i�}1�SV�E�()V'㪱{,,Zܩ[.8F�E��+�@l��(�=J3��L��������"}F�KiR�Bp�vJ��ІO��H	�t^��8H�C
�A�Y-R0e����|�@�E��\1�w�	
c�W�R���~��`������`�y���2�39硃G쑇w�.���*e{�?~�cSk���H�կD�Gw���"{��̯����mϣ��z���|�n?)��������>�1���
�5V������e�:�������O�/,:�w@>��OL7��)�mv�m��T-�{�1��I;r��a����t�^�5��K-���$7zPTp���C�R经��e�����=�����<[�9���m�}K_�re��d�uY�-7�Ɩ�&���m������&�����1[j�K9��˟�\$C�v�؃>ܫ�A��-��ԜW��߻/X���۾u�W���;qrʭ%pU Ua]���X�XTy�)���"J3:XLT�����qZi�܂�:2��`�dn}7X1mk461�p� ()�V\�7����J����к�BM��x�J�����R:x���/O3�FA��6+E(+���N{3��oY��W^�g_��)�df���*�:��C�Ǩb7e�1��
 ާr�c��CV��`-f<[ɕg�6�
�Յ���k��u?~�F�3�{ ���Η���V��}�/�ۺ�B�Fl��v�ȉȔ�U�
B\�v���b�����dT�Ѷz�ӥ�LƐ|����>�����F�e��I����^���UNi;kW<�Z_fG�ǵ�v���~�F���9�m�sX4XV�?�a����A��X_4W%��q�I{##hn&�2�����߽�A�������
��@���:	�em,�����^�:aِ���??��C^��7�´]tA��k�� �`�S�@l	�
�C��7��qA���H���(�B�ě���<(�{��R��|d8(� ؏��a���SRb>Jc�����?��n��\8�(�J�U,E����<�y�.���LA�³�÷�>���r*���&�0��۶^l/���Ju�9���q!��Zf#m�?�On�(���`�K�*V��T����v�R�g|��mlt�6l����똚8�{��ͷ\���ꫮ���"�C�'���͹3b�\j��¿k}�8*�&����{��?������k~��ʾ�m��w\7`��G����#I�t�����
���l��A,86A$gY,-|DiZ.k�J��yN�<<6��I���U���������d=kA	�J��XP�Ƿn��XZ�J��uKД�F ��k��De�G, /��18<�4&R��_�k��)�f1l��L 7͒b�Aq�7���]r��8��ķ����e�(��Q�U��K�}%�Pu 1!Ȩ�`�/:<K/��m[!^�f$�9d�ʒ�1��_���;�3]��& �Eߨ��}�?�Ǐ����g��Ipu)��`OWka�+3G�nt��k��=����l�5�7��-+�ݬ{.�<>OL��ۯ�{������Ïtء����=g;y������I�G�9�!;v�����ĭ(.鞠/��%C�u�����ұJ6��4��[�5�UF*x+/X�,�i��a(ȉ%��R
�-����*2�_�5kW�f&X)��
��9�aSԃ��n�*�����Tc7�蚗=��������4&� �A�PP��5(jkՙ`m�D��&댵�\�X�.��F��J�e}��N�=�¿�c���0K$�TZ#�t�K�{Zl��S\p^uv����d�n5�Q�r�@��g�'K�Y�1̼�pMk���.��r�`���Vm�ӵe�c����50�}�@'=/�����S��?�u.1>��G��j��P�4sQ��I��f� >���ڱ#��Ѓ��[c��68�6"�Yg������{����X���=����Y/��^��0{��ĉS���7�Nǃٺu�kjR�H�"O��*�͡^���ȌtNh�y��M#r~�|Xboy�[���H�� �U��1���
k��M�)<�x|��a�u��bFbN I��,�X�|~|���.@�X���0������ e@!$ș'��
�2߅v +{.��9>� ���M9\T_����W�@V�����C���J�5-�c@l((�c�߷϶���^�ĩ���^��AI�'�
H12*��^ĐY�V�����=�����͆�K�[τx=x�����F�!�c�p�����s��/X�6OTP]C��J�#����z��:�@���l٘�L����p�=�e���C�r�������l'�~E^1x��ȐkV�W�?��a�~���9�m�k9g?��MF&@ڶN�����]'+@�N,!�m���)�,k��+ћ8�ųe�6�eu(��G���7i����N�5�_*���`�Ȳmx����J/L�۰�y~�|e�Ɉm�u�Ќ�M��^N��6��5mө5�{� A^�q�7�<^���C�����\����<&�@��7�f� ��@)��0g�S�
���O�U��b���=�sq�*�3{�{1���"ݼ���k�>lr[��0s�T����g�Ůt1[�*�B�p�{�3���&v"��稩�~p���磔g�~�����>�E�r0�����h�2yj��aϊ|p`8��`?�8<��
�sS���Mr�dYɺa�@[1�փ���j���E�r�������1��Qx��%� iǔ�*��HpG�l��6���w�c{}�S0�cp�K�c;�J&L:9���4����k��a��!V�z�:�8���EN�ų�b��HM��5�����Kҁ��-9�T���lԱ����w��e�h�^_�җz���80�x�"���5��]�g
Ͳ�T�+Д���u�*�4�3����C���H�lWk��y�[�nS��P��b�K��xz�Vu��<n���*�p��u���T:��xN�� �r�ʼ�T���^�y�{�{�.�(��^�w�N�)^)|�Yz ���P'��[���%#�F�sb&-�/fe�N�fy�_�b(o�EΆ�J�5p~�a��}U*8'�PV���uc.|�+5��+�A[�b�M�<n3��
�����T��F����ٯ���K�D8 �`�KR����T ȿE�&����`����վ��3��,��CL@5(	������{�;�5���u�`�°��\`�:7�Tf�F��\�I�~+�o��H��b�9{�A�_�i��[���!�2�T�����#�S/GM
�R�c���m�2h'��AM�u�����}�7�tP��*�3��ꭺ����n�"M&sJɤ���(�L�������}V�>ޅ��� o��B�4�Rʷ��B�"��&�%�M��w�����:�H���q&&��Z
Mͳ�x���݂c��^��ѷ3�g�V�^^�Ƿr�/Y���
_�W�g��r��_�,�aQD �U�+�Y���`}i
�x�u���f�ȏ��.<Y2�87q+���y>G�&s��L�}Z����������x-�̤>~�K�8���ڧ��e���]�:Ԥ�R(+A��	�P
���v�N�H!�L��lN�c�O��{:7= D�!�������E�O���7��_8�D����WK6O��0����yZ}��7��]b8S��X@,l�XNlB�(cH�/�>�g�8�ڝ�X���d��˙k�ͨ4��Ջ�Ƿ|�x1��@(L��Z-�9.�X΂!����W��pf	
�S,��ǎ�m����>���ń��k�����W�5}z�}�Mp��H��~��6^A ��@U��b�]�X��&p>C!��Q'/)��A,�Ua�|�T�(/��N%bX7p;�X��r�t��WD*Z�V��ͨ�ݓ�#6T�g�gڍ�^,+R�g�z��ݷ�H���߽UZּ%�P����t�z�_xB����|"i�����v��t*	_̕�,
����S�8��#v�P,D#�'6���I2O<�y
�,��<��m=�U#��ֿX31��h� B@�����x"|�|��e�� %��Y�+_��(��k�@���Y�{<a��+6!��6�|��VsQ@$�b�s.���!
׈��us}�n�����Ҍs��-K;3��GOZ������И՛���NKy�q_f��ќ��p$U���PBJWr�C��!�o��}��3K|���z�U\Z����Xe����HcbStr��f@���g����]�}�6[�SCT�5��>u�U1����6�)n�~�Db=G�f����0����!�	��u�]��?��?��yV[f��8�)�|:r���g�������:��Fŋ�,9��S`]#�	�-N@��MQbc哵�<$������ �`�������z!c;B�Nk{���hp�?�����;.��1}����=�R�
̺1�윘f��+���b�ǐ�#��Wa1͢��su��q?g����ȫi{č�ajh�*�Gd`��Pڨ�r^�q�[/\3X�O�ɩ��lLY�B5�y&C'�T�f�K����dXv���v�����������3��e�,TQ!���:R� �bS*R���pLΑz��-b7Q���[�kJ{�w�J��G����`G��Ҥŭ��BOEe =~�u��.�0�V'B�@si6;�6u����e60X�L��R����S��~�=��RA�������k�57bY�w�l�'����	�?װ���,��h����قֆ]�*%��!KFCʡ�i�����ڀ9�s�C�Ϯ/^���<�Y]7?f�0�Ώo�L	Q`���N����4ax|�C#ܜ����E�	^��#G���NT��GP7�L9.1+�C1CF|_�\���W���wߝ[�@TdqM�3S9�������A�F�+H=Uj��STM�E��t%��Ub_��`FE^�j^��ʱ~Wῢ_o�K������HcnE'Xd.�ã63W咳��ߙ�H�j��ɫ����N>�؇� Lɍ�?U��-��ۨp��[��0SL^V:̅w��OG��H����O�)O�,����}Ѻk�x� �
�B���Y�D�um�`�5\Ѵ��ULS��� �v���S��Vp$�oz�0���9�$2|=�,�_���9�r*X�_�S����y��A>�&�K �}@�Z�~�&c���d��yۮGq�PO`�� HU%��'q��a���"�H��b��z� �S:���ؗ�={zF2rZ�R?|���޵?Ҡt#����%��2`'NM؇>�1�[+q�r)ҳ��xj70�HNq���8�����kg2�S�]�W�-�ʧOg�*F�`۳^�zV���ز����L�X���l�b�\�X��Y�~]�y&n��CG\H�2m�~�r�����Gg��I�+���f+V(f����>� �o�^8ǅ��Ӷ�SǬ7PX0��N=��<}�X-x�j^㪻���ȩr{�4�$��M�et]�0�|��G�A������w<'�Y��H���� 8��n�B�N˶|�����/��҃8�T��� hUg�⫵���	��ˮ
U�9E^E���[n����҅#��������Kw,踆��ګ���^��<�)pn?CŇ��87^FJO�2>�q�t#́��S�/�#|�68j�����ÐPQ��������V'�g�M��Zu`>�P�j+8w��}�R/8�\��G%�u�!���2��G<@�j�1[Y<�kE)׃bf���E6��l�+J��7��g��/�������lm�-8�7�!�O��v�~}�T(	��8(���]Ps��AҎR�"�Ry�ί�"�Bvn��e���v�ѱ����63q�]ڊpڠ�����v��1�7Z��o!.��OC�~��2t}*����L�I$����jCҴ]�wޙ	^X��)e�T�3p����%Av��AoX���sX�@5�a�"`��w�ݟ�����?T��^���G��H��X�R��<� U ��Dv��Ӵh-�����xq����+����Z9�^.e��ю�9/�(��p��XYO��� F�������U�G��������>+���Ӿ@�(�;�V���W\��Ä�����{<��޻��yH�����Ԟ��:��'�Q�S�*�p�c��\�dd�^������	њ��K����6�zԖ���۷�'?���O�J�E�+���,���jv&�h�������~�� F��ќsvy�x���#v|�DX(4np��J����-"aQ�pN8��eC�Ñ�/���,n�w~<�!.~�������� G=��D�),�!/(��5��Y���<DV���])"Y�b��wxM���f��*૶�i���֑��hX�Bܣ[�;y�n-�:�Pj�~�]s�e��m�;
�v���ܲek�˷#)�"B1#���6��R��ѭr�s��
��`+3Ii���]��ee�n��Y�������;^���	�j4Ȣ[�n�]{�u��ؾ��/�}��i���a�I���^�{D��۞�^�^Y\���ӮZ�?3;ִ=t؎�<�^��Uk���>P# �����0H��{���ܕ�7X��>��O{���:�&���`��Z��ێa,��R��������U�"�x'+Z���w� �W��I.�b"K-��z�<e�S���^N�x^��d�H����~��7k�կ~�c�<?�J��@a�b�s^�5�)PSz֥:�!�H�T�#�X ����Z���Utυ,.E@�F���9׀' ,�aD��9�3V��?�)�Mk�i�,CZ�Qw�(f����Ms���l�����٘v��z��s��@�o�{,��(OJ��w-S������x�N瀋��	o�>�Т�
^��V�U\�ƾ��_��_��m0����U�7sYr���z����.��U�9v�O�S'�z���������}�P 2<4jW^y��t�-62�<�Ղ=�Y��Ŋ++���@Ѝ�����@�
�Op�~}���h�z�С����o�ӥz�A�"��l�s��^���^@7���\�;��3�"DbKq?��lY{jB�TF��.E����xr��M��`�eRk{��g�D	M��q8���{�oe舁�2(�3����Ӆ;B
c��Y�<w�8�a�C���j_P�b�NF� �C���"@�F
�O<asF��c��I����7�r�l�!Q�_��p��o���N���Vl��Q+6P�ᆗU�
h��Uʶ�.{�*k�>�2��̝���E����a�L��=�;�p�a�^{������g�|����m;l����-ۂ2\m������c�֌�ٛg����Ӈ��z�_����ş?��˯�ʞq�Mv��^���G�O���/�q�gT�6�d'�����^��9��%�@)da��*'X�����������{(ɮ�\x�[�s����F3#�r@�H��g�c��f9��᷍��l�1^^��<�m9'EF9k�&O��t��|���s�ۧk���i�3u��=]U7�{Ύ��6�<����je���Mo���IY�Rs�̝�d͊3L�U��et�������?�	xu1Sis Kt����o���`�ca�} 3ȹBW�
�=?�%�aB_�(���H�Q�.J���C"B�j@��ר0� A�
���8����y��F
! ��~���8g2?���*��_+}q]8<R�EeP0`�1��4X�^�O�Z ��������Bޜ\���n��f�sޠB�O-�N#tC���4��L�RN8�@�2U7b8�f!N8-�\G�n�e���O�s�(;�C�w0�Z{ը&O=��<��C�k�.��^�z@
ټK#r�����]���x�,Y�'���Q�������cn<Щ/��z�����JcґO�����X���e|b�P4�5K�Y�bqT���?��O��x���C��&�Nc��R��8L��$�Fֱk��X��C�����=%�܀���C��<��~�;9�6�ɪ%G�`4�^,�-@lѕ�H�
g
v'�5���k������=7�	�P1���;`�d!a���I��*]��� ���� � X��
�TL��H����9�]<�&X�P$x���964�EL����E�Dx��H 7���Nd,�b�sa����f��`դ�W�y�j�G����Xo{:�^'}�+͍���l\�Z�5V����`�5,6�D5�>�A�HO�ׅ(����6��R�A��1��wE��j�T+#�����HWg�Tj�תқM�T�.G����?�o򋷾NV�� �V�4E�o߷�Y�/£�4������4�X2`M���әH|�ټI'z�2ٻ���.�0g� d�'&�TQDr�h�/49�%,X���〛qO,v4u�{���bs���l� �U�������\WW��s]R�M��A�KJ�c�D8�U�E
n��K�5
8�t� ���%*��%� �c��AE�nPldN`C7��P�q~���a�@���j@b�x6pg��W<8'�)�>1�sM�"�����H$*$|��̑����)�	�m�b�i�G^S��Ϫ�*�CU��Ra�,{x��}Kep`��������S*X��Bz#n����Z+Y̽\.�1\�=z�GO ����U��ɸn|�P�z�>���^�v�^GE&ը�zGw��G��d�X�cE�_��l���39s�F��{���q-�)/�-�6��BQ+�V�IOW�.��F��$��QT+n�Z����,��`��,-kzՄ!����P:q�:��Z�܍ՔH����w�i�6�&Zp�4'�[J�$"��jm*!��u����ez�hm�|,a��.X��Wb����,m5�^ ������sI�8�/x��$�&�V3>%�����B4�����}�vZ�Q�!��i���W,�����J�|�FXc^ ����������a(�C�^=6��v|� �C�^j��](��ߧ7�VZ��Ĥ|�d�����T��	|��޺�e+�������·�#�x1w0���IÍgxp�n��s�:�3���ۗx�&9
������y�]�s���M�����c�V�ϼ��Z�S_��3�< &���C����
�:�L6�`�@b�V�,Zj�<>�)��vx����}���l������©N[s��UX�P�\-
�x�FT�D0
x:���E��~*0�7��ix�e��!Y,~��7(YI�CқL�m�ϳ;��v p��b!+�ɷ��h,�:E��!Zm��S��}�����>R�gx\��a ���&�}( �����8��7�zQ��(�ώv��U%1X��~�a{���G 
��f�}	�j��`�խ�5�=��-�S�խiz�܂��
����rV��� k^@���?�cy�[�j�-6�G.�=(?��֮6��e8�
:�!
J.�1T!
��+�*Γ���Ge��{�
��x)����@��#)W���V���|.)�w�>��^�x`���QmG��.'����Q�X9ࡀ��ݿ�8���˧��8>��J"[�#��ȡ]r����EK��j��Er
��"RQ��"�T�z��p�� ��A����	D�A��ˎ�c���T���2�7x>��b<|�B����]�Uxn�,~"�$�'����r�}?Nx����Yx�n�v�f  �K����
}	��N!\#'z�8P>���:������nB����?C��D�W*��K��uOEe��2���C��t�%|����6�~$�VUϿZ	�=��S��;�}�{���pohbO����"e�'=8���f;���T���CϛM �$��>�1'�*�(F�FOθ�f1���9�S^��4s��ɴn�j��X��8��o&r\aUh��x�u]p��@�,����x��K�\p@䰘QJ�67-Y=����=\5i�8�o�^ߤdԺ��"g��8H�X}GӖ�v�K`���0g1�5v\�\�>�*?XC��;=dȇ������=IZ�P\|nx�a�@��eX��C�/��&(4d�� � ���%+������u�p�����Q�Qt�B�v֔�|w�}��
��q���ճ���o��8��)����Uu	t�E"jm�z_wv�˹[/�J��*�T���O��_�.)���@٤Ru?���½c�c[%naZ~���?�01o].�V��~	5��ať*R*oV�[#Se��Z/����i��~�m�w�AV7+~���~�*[�H���'�L�w�v�Ly)tvYy�Χ��2v��i�+҈��G������w�y���w��][����f� !� �a��tv�?2�o�BKf�4�Ua��EO��?��B\x8����Z����`����2QeT�~�C>�>�n��,ߘr�J�g���b�����Ig@4
�:�g�BKPX�;P�q����hL��a�T�����60M�F�9i�wS��EE �z&e�8�9���U'`1���H�m=2�����,�G  ȥ ��#���!�t�2Y�j��Ke5�ft�ܪ��7�vmM���5�\��A�H��}�z !^.��������X��v���-MUd��{e�sd|�\x����'d|�l�7����V������(H\��7�� ����E ��<������q`M����z�굌��ş�2z��1�4T�hp]�J.Hjűw�q�.o6\u�<|�zX�،p����I\��'6:��yv����ρ
�O��sD��B���0D����������v[�x�X,#�^*��|����W��(8*&�휺�p����w��@���>�)�V(BDØ�g�ٱږl��
���˩�V��=�#vC�����C���0%z(#B��q���l+a��6{`I�Ž!���G>��%�5p�}�c�R��m�](���P�ꀾ� �Ī�e�Y��[&�;�-�$j	�=���
��?�8����s���A6�K�bz?�C���iY�f����*��2tx���&&F�d,�.Hhn�z��u��$<?b�L�b��� ��͞������&]w, +��?�����~N]��y�.�$��8Ir��K�\i�yZCjX�ӷ1/�5�����p�c�(6g5j;����$.��a�ǯ�3���%a>O˟�B�,c�8�6"餱|��iE`�g
��(?���{���!A���Y?�����-�F/�`���U}�X=�%r�Tn�}p�O�Tq����L�#\w�QC�� �_��_J��0ҡ�$l֧� 4��u���Kj��a��AȝBΘ�׆36�5��h�ò����C�䓻��-���Fr�q���uq��>�e3/�FY��? _����u��U�rM]���iG<p׮r��ak�GͰ^��Ns)�q�C��p<��|�3�7�Ɋd �#�V�+^�
��W�l^+�i]�ӗO�v|R'��dCv=�CjU��֝��@>+�5���E-�T:�����Xp+�%��'(F�W�p�P���'��yQ��µ6����0"�Ճ9gXe����e2lCd�X��7C/[�Z�:��q|&*B;1��҇g�d-�E ���Bx#�okk�81i��By��l��R@�*Ž�F�#m\�į �݃Ec#�q���ڄd<�1�E:e׳~
4϶XQ��������A��0�BD(��Ї>��ϸ�gp�DZ]�{�!�6�����J]��d��@�����<8j�����l�v�z,��� %�m�}�d��5�i(x�q��V#p�bb�(����N)td�%/y��k9Ier�eW�Y��&IN6��*�U�����1w�?�c8tP����ֹ���k���H�R�����k������X��Q���]ۤ�_j�Ѓw�#�X*�:�gƅ��J@%�d�.�?�.�@�a�<����r���ܡ��pNl �5躓��վ�L����7��S����?���~׬Z]S�@y& Q�=6z̅�j�%䦳7ʅl3c�;`�j(�񊅐�� &�>rԎ�Y�0�rd�����{l=�
7(�8��EBki��a����V����P 𤡸 ��}�8�����Xƫ�Є�f��ի��[��FR>�����è��F�[^�R�3%5�r�K�������ռ�`<��/���y9�c�~�<����84��+��I.[-����\�(�~��!�c`rtJ>����C�<x\�x�(l���s�J���}�0�x0�L���p��T&�~��񉒹��t`�@�����pb�@� ɋ��x<,�~c��*!��.#,�|v&_���6���ŴI7hd! @��
S
�C���,,*�zc���D�c���  �ň\Y+`�!,�{D����m�/n�ه�an���<��>{H�;M�	�i�3��:,rҋ�w�e��_�m�ug�  q���7|���Hр�`]�<�'�>�{"�k�9(!��\ӣ���v`|8+W,�m�oAה��!�`�aF&U�wu�[���j7xwu0���$���ɸ�g쇛~��O~��	����J���M@�Q �	��,�[�J���$U,tv�cO<n��@A��!_0׋Aӝ��?��e؇}E��"��K�я~Ԅ?�
؜�dY��H� Ə���b3zǬ>,�?��?�ςW�f�|�4��bq�����gB��⛵:�B�T�'Tk	-��h�`Ψ�Q��m��CH���j���.�s/ ,0Z��� H�`�ạ�|b7Ɗ�����i|ZgZ�0&��� 7���7�O饢0	��[�����ǏkA��A��w�wm���_��	i6H��>��4��:X5�A�c���뿶�!��ϡ�PQ;T���&[�c���9���i�5b�sd^���p*�^�Z������\���s��z�"�^�|Y�|�]���S���j�Q����|����8��q����D����d��/����b��)/��d#$d.2�Ҙ`,>L>�U0�c��7,J��ȊȒo�ƳM#�}>�O��C�~��`�����;?��D]E��=$��b�r�@#�nD�"����C��Q5��mm9���h%B�����_h����{��d
d��j���XD^��/��`g)���>�|����h���a�\ ��{�]���a,����`������8'�C�<�������ll�C>�=7�R�,�FՅ�@��ϲ�{�T�޾���⹌�=��F	��� �R�*ܔz���?���9E�0����������=<G(W��^ �'�7�1�02�9������:��|�5~r��˰i�4�7��eec���Y���������0��I��k0�E�&�	�釞����EuH�<��s��0���Ca�L���U��2��m�ԋ��&|��ZG�o������m����Hos�~��o�+��aeb�A�����p,��/�.,�w��]	���!�������c���#$�Bˇz�ӦWɦG����i���<����M���Y=�U�@���7��ֿg���۴Y���K��[R���*�S���64�JK-UK���~��Y�HH�sG�������C���O����-���bIVi3�@�EzrW ��S^��7�Z�/Fg��������d�9��O���,6,�>�$P��d �Gr�%����o��L��:J�;��뒎�ZS�qݼ�p�k�}#���:�7��!��	��[�J ���Φ����>.��8�AC�\�X#C2n����7���a"EaϺV���%��3Ɍc5�c��B�'`�1@t�F�*����A�ǳR����'���w�Q��f?3�Dm�r��V�4�����m�:�+ӎ�>�0}d���������w[��Ph��½HXã�L���C��DC
���3f(��c���c��b�i/�1�L\{̰�9>���
�Ho��\�x�X�
��P ���U���[� V5?ϟ�l��l}���oTC)N�%�B��KnNʕI��fBG�4R�ؑ�ſӨ��F����n��D-�b!j��LaDWߧh�����rV���X}�(r�P �*��q\*,����J���P��	M�@������@1�G\��J��%��ҟ�]7Ce� <�??�R肇�ew��fA��y�汦,\j�9�_��P��q��=�1�"(?�opݸ�}�c���7�5��"�3�O���lY$��>�~=A+l�?N_��<��R�\Z�\d~۷Z���9c�<-��H�!��W.x,j|�)3�˦|�87,�Z�YS�	� ��e�?��q�wa'�L�l���j(�0� �AT!�,F�i9?l��>e,�n?&;�:k��(��!�?��}( h�0�DCk�	��6\��!b�T4P��nR�!1��3�l��ռG�Q��8��CD>�r����Hv�V���!��c�L�d��P8a���֫�7���q�?�9~��=����?��$J���L`ؓρ�<�$������<��fΆ������Nߘ�|�_�>'6�o��	�kCDxDJPX�'j  �a ���[@̵i�$�oq̮�&�՛����~�)�nE
9wO�c��6E��[D���,��FvōG+�����s��%�[t�3n���R{,l�����/���6��/0(�0����g���}�LBC�x��|H?��?�Z�~�����ѐ	F�/s]��ܵ.\�а��Z��n�\V�"0@�{F�����2�t�q�)��2K��h�^)ǐ�ؓͪ�E�\<Yw]4����	��g��)�i(����7&������':N{����;���VN�oՐۃ
�V�����	��l��e�p� I?"�=�S��Q� ��PO���ftb�^�D�T���F����9c���;�q2G�e��o�QPxFC̅w�1��\���;(MT�T��F���#�?$�HoϠ�^�A�U5�O(N��%��f��	z�T�����"bh�ъ��|N�"�@Z�E���IfB&9�,�ހ��i��!Z/P���s����T*�w�voeA7����r��n]��DTܗ���V��Cf�l����� �Q7��@7�Q6��+Z~�M{<W��kQ-q���ټL�F����K��ua�Fv���9cI^�74tHB$��h�3�O�"�3iT��4ʡ�-�8��a蘈?�C3ĕ��Ӝ�8��|��ӧn�`�#Q+��LK����f��|r�3yǇ��{<�}����ύ�$�,����T&[z�r�H9��(t��
c��b@Ӏ|�]}�cm��8�cv#��]����n���o88rW�Z:���V�e]]0ҜYŔ�4 %p�l���}�*x��"F߈�	^�b�:��̣�8i���"=�٨���4����  ޘ-.��Td8�w�h��°-v��|<.CA�|~a?��\�KK�_�R�ԪGb\+Y �b��Ѐ�Ti��LUʒ�,>ZE�_��u� �'���Ӷ���6f�I��v�t���)[S&4a�u>U�X�s���|Q[H��ܴ�vh��˷�����'8� �a�Ic�0�I �oȠtj�{��TP �L�_?Q�[��<O'2Ny�?''r<U���3���	.�����Xt�(�}aތv���Wr0���#�J�xD��k�f\%��
�TC,�+99U�kba������7Bc\�f��Ԙl&������h��5Z�HrhX�rprj�5H䆇G��Iވ���d�*Z.�^�W\_$v��'KR����d&�l͠��p�&�g�f�0����~Q��_X���F���?�8��f��%N�D
pChd�3�A�؊�������a�M<N
O�]��Dt��&u����bh)���D[��{��T,�F(�uߨ98_�~�]����I4��26Q�#G'��k��ϿVV�X�\/��M��'{�Ʊ1�T��w:�����ό�J��zcK]��K�O�I�Z3�P+�Z�
��:T�ҥY�'P�����U2Ĝ+:K��x���]�`}�^����V�Npq�fU��F�m˿����� T��1�6�\�p��er��73X��&�7M����y��կqpb��)Q�ҝcl��u�`Xv�6�Å!:ؔ��y����ʰD�8��1��;��T2k��U��C����%/�ŘH��5��7�~'�W�q<܁Mb���dE��>�d!�	��A�h��Ȯ��Lޗ��I1P�g�t�������6湟�;��u����毙�ol�56wMM�y�Ӵ���<���6&*����<�Y�ef/^����Le�4,z��Ҥ|���_��~/e��W�6?�/��[�o�Z1A福u?�@��1�f(�����8P��`�.�#�����d�gZ!�o�:����ϒ+.�\���oX%1��(�:����x�Є�iZ] ������U����'�z����1{9�r �=}�d`�Y��=�׼V�{�L	�(+��u�Ԫ�U���#�
�Ը�FG��L�wMi�Fdx��f#2%e���;W�V��b���d�X��K�����G��^3���
�f:���2��%�Gk@@4*��<���(x;���T��3�!�V�7{���ǧ�f3�ڨV�,�0��,��V�..�!"q>���n�.m>%g^Ohg�3FH�7�����$��$�%J�e�&��I��H�V^q򨤲*X¼Y��;0��E�S.H�����y�����y�E�P�J�)r�/Z���@��@?�D=Bz@�`/�3�Z�l\n&�c�PF?�FG9mI}�&�׆�J@�����u��<Fz��?�����"_E�������Ƌ��c J�JY3p��L��z,E��V�?,GF�4b��.3�4�'��(X����Z���L[��D������7��g2Xc�$��|�͇tC	ԬaRl��=i^X3���X�˰k!�]������(��aPV6tx�>�d�R��R��Ȧ�Ζ�k�[�� ��ߡ1�N�E��E^QԂ��r�
\;����*��ꄏZ��O���k�����I���/�X�ٲU��XeM���j�`e� �h�fO,�׽�u��YD���ˇM��D��d�"����0b�ȬE�o�,��}��45i:������czh>��kL�h�!�'%&TL(�@d�d:�_u�?2��@������4Bm���7��u��b�/�G7r���w�h/��y����HP��JkB�}&��#'\U���&�èG@��g2ܚm4 �.���\�}P3u`-��}���~?��*��ç�-���	BrhP
�j�|̏��X�7l��Q�h��dVn΄P�2���Ϫ������ร�_��-�E�Е+_M�=�x��GT���8~E�F�u0.�鄷	^���GS�h�X�O+Q*��8�c��T��p����}g�/���(�}�1t�1�U����T'z0'&N����ȇE�?�}��(䬝㱣#*�'�|\�������q�9r�ŗ��3j����?޾=!������u:7po阡�I� [��u�\�|��pJr�H���%w��=����K�汪�h�����^����L}@Xl7�|�qsӊ�5 �>r�B�;���<����_�z����[,c�� oj�+����Mق���"I�b¬h4��E����&������|�=��A��t#����ZY��U�(̙�`a3��1��V]qI�zL��n8P��YG��7h՗a�=4�?	��x�e���sq3�,��~���5,����F�	�Oڊ�,~��±��	Ⱖ�جi"OƦ/tmQ���҈��A6gE;
�nK����������R��G�� U�j���5m�tʅ$Cԩ��~=����P�t��$���g�W�<AJ�����v���,O^#�a���$�3��E�Y�<f��;N83��0%Qz����Y�C���k�5FS�����@oP���������߃�����7!{�<!�|ر�I+P��p�9,O��>����] ��Ke͚U�8��'w<������I�)/�[�}�[M��<O7�9��f�c�%���[�˭��"F8:<l�����_Z���{�g�a���2��6l��.���P�o����Qs�����o���a���d%8O���>� ��:�ıZ`Q�*�'�N�B�gI�,�����QF�$�Z��W��I��.����P�V���<��*��n�JY��B��9"ׂ̡�G+�!�{� �Z��j2�|H�S�:�[��j}DJ�q��(�5e���;oT��Vc�!��]X�8_Ը�(;u�"�%�!�jჷV�U��KO�R����E�*m��N��`mG�0�9*�ָ�U^�q�:�*@Gꗊ��Gus#�l�r΀���V%�����U3�d�ff
�|>Ãa��-�Vፐ_:t�j�ٺ9NVV��6���
��e�u��ީVc~��ǯWFr-�����Y��>��"��L�����`���"��_��������@��=����j܌���!��I]�����3��(�՛�*���-�7��笁;d���0W��
~�S^�����q�s&��͛�ڄ���ʷ��e�ֳ�uk����	�6fdl|B����	�y�u�]g� x�Gy$�h�F̎�V�h,�p��2f�����2�(�}S*�U�,D"�j�J�B4�=I�f�E+{���M��5 �j:���F�4�.<�r���g�/��Jy��+׮P!1�B<vC�p^�:@���ty�*���q����խ���C~�
��� E{��321Z6�epi���,Q-���+��v=.���p�K�8�B;+K���a�H��UUL��0p���T,)it˝j�g����#�^�#�s�'���/�;������REcޢ�wthJ���άtvAY�1<�I��g6�#E}��[��u�ͥ��)�� ϰ&��f&k��,��nTu9z����O�9<t����N��~,������cR���r>��I{,�1`U}cF�k_l����8b.�Ǽ�����n�[ �B���z�{�k�;�������=�\�T����񈮑��Y�D��)kh?Uv��K��������;�'+V���/���m�'���>�ih�e�<兿��� ���U�;�Q�������q:\(&�l-�p��B�S-�1k�v�-��%�Nm�����	�^ U��݋�/��/��@7%߭$wG3�ۉ�f:�f��E��I�m�ΕMg�։�������*�.�_7�V��@U��C�F�;������b�'��R#�.�ۈ�#uRy+V{��G��w���뮽J��ҮQ7�5��Z�D�#�������wn����u�Y�e�:U&�di����*��>V�o�^��(ʍ�]%}��t�۰�W#���kBqa�'Z&Ǝɒ%r��W�v^ ���\�>�HY�ꍤ��Bjt����#�ߴ������*.T���W���[=� �8�s5>V�o|�G��^p��?�i�/��!��IC�c�׳����m�,W^u���Y�9���	�F��R1���}Xʓr��[d��:?u����[�}ʱ��7��GF�^���K����<��E�����0���V��O2|�B�������~�+v.th����Д �������#r9C�航���xTe�r�?��q:R��2/}�K���蓣:Gw��r�%W�~h�ʕ�������f$���k1Ny�ߒ�'r�-Xh��Uj�8p�ڿ�P��֩��::T"n��*�qO
ZZ"����H%
��;�y�?��/ؿ	�d���\�6�
�|/c�O3���#maX)(�)�&�,*��zք�6>Si | lr����VQ��ch��k��"��Q�o���@Za������MB�%��e�S1���ʢ�	ز*�@/���`��-��p�f�︡�
�M)XE����q��B!{p���Y�5w��]C e@��oOA����Gz�s"��a�,C�j��u�A��~�
���B��Tծ6�BөF$��6�8!�Qu�"2�IxO�������Kh�fG��(���e3h2��zQY��	bNcsGx����p�0����@	�z���Hf��q��b�q3RH���kD������F$�eMJ6������L( �u���
�9��!t!C�^�7 �@����/����jҮbxl|D��R}�i[��a��	�$��󙔮�kk�DgGo���:�q����o;�����Y��h��8D���ߑ�!>��x8��@1��o�����P2l���|/����Ic4[K��ɒd�ŵk�yF9�؂��'"5WSV6m(���+"6mEh%�w ��<F�v�C@�@�{�X]��Z��[,��>+��Q$�1��	,$N+�)��ͨ�"1�#�آ�N@:�G�a��į��\�ؘ�rQ�6*��UХ$��}�*$�E*v�Z�b�]U,���M�EU�����nT$V 4K����ҁU7!�S��͍����`���K��T�~�
�|���ME�Y�Q�nM|`������*�lƞc��C��)�C�-}h�':ȕJS�iK�?_���3H�\�F�"�i�0��.Yh{*c���ײ�D�I�;K�B'��b�'
}�A`�{�{����ޒ��?��^�*���lﳾ�͎X=��Z2��^!��kA-i�$���&��,��`^\�:��n�2��3P�Tͪ&�R)���>�.�	F��	���v+�5	:eCnQb��+-g%=<�^z������7-.�������/}�K���`˾���}�9Z:���9�9Z)��,�kp/q�˨��E��*��:W�Ѕ�`� �Ě���3b��#��Аad �g"V["^\6��x,���5�Q�)�@b��0F��s�H��0��$���g�TW��6��nө72U���В�����d�D���x��A�ϪL��.�	(�sʚ�l?D筼���E�(��'	q�!Y=^�����2錛�c*劕j��	{�~Y�5m	_�S�u��z�����\C)�)���=8�qEP�_#w�$�[�<s-�~�O��a�Cj��:m�P�r�����Fw�>!�Hp߰�Br�gfM��c�Ν������oΫ����q���8�RdH�l��F�*U5�
�NWcr``�<f����=.'�E?����?�@U`GgA�����Kz�j���V�[�{���Y#���L��DE��V����6����^ ,�������K��+���|�#����\@$��U�ܠz�6}͌��۳5��������B�)uOIU���`�Y*X�CG�&�!���F"��F�j9v���\�g �[�`�a�NQ֡�fE̽��N����D�����>��g��ʆH*������g����1�u�������]����%a������5�Vv���W��UG��r�p��BcYU�cG�z�D/�`�����16Z���^��;t�����|%e-���hk�3��8����
Wmj�Gz�X��$�#g)�JU+�����̑#Cv{� B38�SQ������U��l~�z-׀�9S^z�\u�T&&;,��/��B������wK?��Sjh��W�hG�L�2#'��ǖ�+����q��gn=�Ċ�0�^��D w��;��p��� ��?k�~���uk7ȡ�g���V�����n���~����I)�|��[^���zpL'ͫX�8�$�%aN��54я�s�v��7�+�-W_�y��{���.��]�K,|�u�u�M[Wv�aX�F�W낯�ӟ����P7�t���o���0�~s�"7�$�o��o���E鉺-� p���b���˖���:Y�|�)��v>)�?-S��%E��EY+r��`�2Y�~��%�?�^FT��ԣ���c,�L�
�^������;e��5�v��1cC>�o�ZS%#��d:,�X�5 �*��'�fQ-[�Tϻ֊���{Z���%�)�\R9C� {_l7��8,��@��߰BV�Z/�� ���'ǆ����,T�kjD����������2A�D歹�T �-Y�v>*��~R�"ٲ%�%U�L>�)� B�%�ӻB֯9[ϻN��1����U>�T����K>�ڂ�)���\��Ⱥ���Ы����?�C�ј���p���R4�����}:��e�ʵ����d����Ԩ	�P�	sVL('t��Pa?�B�]+T���9����^��\6{MHDW��؈��4k�DӍ��j�}�8��1�.��ϱc�~��_��_���E�@����Rٹ�aٷ��Շt��V+��;��e��~y��'u�����,�F��@~ͼQim�EQx��}��#
m��bR�㮻�˥_&�j�#q�~�9rdhL���'�ʭ�1n�p�W˦�ےb�{��\>Ұ����`�����|�k_��Sf��1��s5��q�-�GN|D�C=!6�I�Z�Thde�곥�g�
�N�9��aCڬ��#G��sm�����L�����9c�f�����W�궚
c��Cf����X��D��2��@ϹV֮ۨ�YH�3Ղ�{߯
V��%��q�����w��sW��X-����JU��U9��rŹ�, ��^��N���M�.TA![P�Vz�d�؈^g�u���oZYU+W�wْ�r��3�"�ϓ�*��� @�*F��Qv�O*g�w����z7���*A���;/��R�Z������Wb�@1V��~�w�Z�)Y��G�?'?�~�
"�ʺ�v�zC׬�?��/���v�U��4 1ͫE�~c�����x<nq��-8�A� }Fh�۷\�:{�z =�,;{d�*���wD�1m��P�5Pn4�T��I����ǯ�hQ+Xf���]�z�z���~�����Χ���5�y�����}�3 ��[���!� $���սT���(���W	dr��Tv��~�U��s�7�h�Ȱ
�$\dJ��1:s�Q�Mҭ��#�������E/ԍ���^)W\q�Z~=�l���[�����.6K�/~�f���H�7��|�r�ԧ>eP:|�w~�w���a[��,�&�n!h.6���.���A�U�ꆯ��4fbq�n������.��YQV�ZŹ��~��4\��b��,��IIO�r�n�ֈɺ ��(O��c!�jC�Z�pܜ�TEܻ_��B-�^�2��M�b�UƻU��ˤ����T������Wk+��2���:u�;:���c&�sªY��l�*1�x����kM�@L��V]�� ����4mJ�����0�TC�W��֯�"#c���ڛD�4��F̀M���):O%��"�*�^�R\����H�`���z�=�dD�j�58�ӈg;Σ�s��J��Y��jYv�K�=�d�>��S%QO�1�U�T�w}E.o��z���Md�h�=�R�3�@�!��3:��~���X�L�
�Azy��y��F��Ac���%�F��<�P"�x��<�b�WR��q��Ss�2,tp}϶��ׂ�IՀC�����?���z��PBr�礝��<~Ȋ׼���[��,]��y���}�?�Ò����r�5�ɖsϓ��X���>�_�)����e�����?j%�<��U�� G�O"����)/��Fc�V���kn0aE�Sk'�ﰅ`t�z� �	d�X�@�� �9T��;��~�#y���-+W��!@iU,􁲦�O�2>Y_��X��<��,�zF^���e_'�ͤU�Bh�^��
��7�u����׾c������j��q�*���U2e�6�I�KRQ����m��yz�nٳg�\r�r����E��`�U`���{���&J�Id�����˱�1y�^��?_�EQ�mJ��
�@�W��MDQά�~���^��]�����ea�[o�U�٣Ϸd��(*������yq��n9g�6����S;���[/���&Y�r�Z��l��.[c��)��`�U��7�\6o�P��|�;ߖ��k����s6� �2B2��&�`EYl��h�֨�c�paC��?���ۥ�җ�D��id�t�B����*r5j��]{�z]c��#����9�\ 7��")輢�"�Ϲϫ�����R]��.ٲ�K�~�K_�b��oy�іXD�i��_��z��]��D�r	�^Bk�C?�ӞY��î}&@�R ,�\�
}�pѡ�:��S����ȵE��>X`����@fpO���� Q���A��k��P���s�̳Αo�9�������iN��d�$w�u��w�vɫq�~�1��g�o��=MNy�H+Ӡ�����y)����|�2Zg�;� �����N��z��g�����.��� ��g�/$w�	�C�ŀ�x�Ï>��lC�a,Z�-��8��%��	�@����Y#֟c��� �DW�j9��F������r>2<)˗ʹ[/�u�W� ,��ZX�g���Q��t�jA����19phH��v�
��,TS�ؽ
�2b��4�,H��D5�9����e�X��.�B�ظV��}��rV��87��0��eЩ2��Uo�wTWJ�l��X��b �ƘP:��0|Y��2}�y��'Գ�+�ܢ�|�����Vv=�A�!��"Jg����S�6WeAP6��@t��X�X(-g�EC(�]w�t� -�>�J����BY��K�QŠ�H2#4�0�Td��U�۷B��T{r���?d��\v��5�B���<G�0���e��Y�"/G����[^�U6��Y�*�.�Y�8�"��!��ݳD�Z�z+Crtx��vδyH�a�#w���q�.V�������9�p�ؓd�D�Ίeˍ��!_|�W0 �
�0��rYX���W\j�H��;�����s��##���ʑo盦T��;t�M�1WP˜^��K�<�pp������Mem~��ߕG}��;V�Yia��jo�;'���wВ�۷ߗ^r{�!0v��8>��Z%0*{�0�)|�S�4�Pr瓆�ս�	o��<���j���f�	*#n�r	N��']B�^u�!�9���㐁�$2N]-�RmqC�����@,�6�Ej�Ud�h+��JĪw+�X!mU�)K�A0cn�F;²�LNLY���c��ڋ�W����jgü�[��l�f��A�r��>���9���}��҃Ŗ
�"oČ��Ɋ	U��1cNZ�8�\6o���*5�r&x�:�]�H#�� �',i��@11��h��C�P!]��˲���c�5㺪��X>��Ƚ�T� }�g4:6ay�FX����n(��Q���x��F07C��y��F�,�B��R��ks�deGGg�9|�L~(R��=:iV�Ɛ�(YL������>"�"�P��8�~�Ϳjt ���� �9�����Y�c�+�
|�+_��M�e��.Dɶ�!Tv�ܽ��ͷ�q��ۿ�h��ET*1P�1�ZgA�����.�
���"&��V t��
�q��׿f�<�:� �U����x����ZR�0��i�� Uox������k֭�߻ݒ>��� �/��/m��B�G�����E<F��b�%����͊�@�WtE7i��8��u��L�"���$q²��nk�ё�!�mxR;G�GIP���0�՚��;��B](	�x�{n}"ǜ�U�?.	Cᙕ�QRp���¸f�Op^��
N��������g�{�.�7N�ȑU�K7�y+�r��(�M�TP�������I�0ra���Ūa]���)?\c*��Z��t�
�i�hV��P˭jJ7g�s�X�*�1Q��-����F��rE]��F��%��I$K5tךN�cZr��A �2����m�y_4��i����Z��>L�r?��e@=�?~ߟ�
X7d�>�Ʒ�������>A`㻀h�3�l��`�=�z]�o4��5BX00-�{�-	�#g\�l�m�>�[��X��c�R?RO,k��uu��B��[�(�B��׿�����`0"��'4>ڴ�9��2��2�4����a���&�1�npΨ� 4��̊h#$R��>.�g2nz��������n.X_��������/����!��^ ��@k�����2I�)�K$�`(���>��D">����2τ���["�P�g�OX��ݜ�*DQҎtnn)Zˁ	m�1 �,����"b6�~^㣅���ʙ�U�m��3�<S>������ߟ�� ���>�9�� ���D�^Ƴd�ܽ#�����T8'�|8h���s��6��aʹˎ!�3��Ȋ���ݴX	�B> E]�Ї�w����躄M'pY��\W���~�17]�t�O{ܪ�Y84�No|&:_���{Z��k��5$>����54�H�s��b�3���b�}2�{籉�'j�J���G�h���量>�-��AZp&�G�b�mmb�B�`O=�>��>�k����}�'��Z�v�F�욟04��W's�s�<�,��:�+rv�x ��>�,9�0|zOT4Xg8����|��8�k>�|�M��40��P���zh�aa�+`����O��L�=Sc�{&i-S�(Y��s�P8aP���rS(���>-5�"�{���M���~��;�w)l}�#T���y|AO��S���Ӓ'j������ p��2!Tدi~�|^�5�3�p[H�p<�ab��B��ÿ���.�G>������yoD�  b���-/ �
^��,����Ƃ� ��c����hNFs,�����ɤ7�'�m�i�yc�Vڇ?�a����}�����͍�>������7�s���P��L!�6�/�}�I���'��Mkʷ�\«��"6Z��5҂Ǳ���hnxc��y_�ӛ�s$�Wz$ �W����d(�a)���򇉀�����2���sH͖�o����}�~Z$H�4?,⯋VU긎�DyF~�g���-'k�f��u�w��N^��#��yDU?��y��ו�W�>���4p���q����O�
�h�%��Z9=c��
[�M<<�������>p�xA�#�e�^ ��6|Z�'{���!����+Z0��Z}��D�-�wz�x�gU�|�<���r��js�z|���|___b�3�G�L�B��p���A9Vw����������\�����4�3ŵ���yzE�Z����q�B�
�G����g���O:8�4p0'�(j��Q���ż�Y��+Þ�������9�=��Z�4<V��6�ۉ@�hٙ���Xsq/��/f��_d�6`% �	�I<
��M�\�}ف*e
!*1ߺa��0U4� �.9|d(&�j�X�͞�h���	�5�����c�3���5�y����=2|Ԅ�/����A�{�@b_���{�6L76�o��:g���Ő_�`}߁�"�s�u�b뉰�ߙ��@@�Ч���5%Z����>�(]�������-,��c226*ݽ=��:p�����87���8�x�~���:������>�~�]Ιڢ�c��:��,����Q"�S��[��g�dz���a��k��c��h�y��j��Kn$n�<^�uIRaa�c0AI4r���'�]��� �}�In��7�Ip�����l$b����L�����hY�@K���b��ap�O~�3�r4�f�Oa���.U�B��U���3ă�
!��.`�Y�CagB ���x0����܎�s��)�}t�����ߏ�7���00�Al߾݊S�5@1c#oT��n�5����2����s�d3��*w>_*zz����yP���<=��Ѝ�Ȍ��}���h�Od������ډ��L�Ml��+�u˗��Ń��H��p6)�
y�)q^�8�no��	&?]|�~8p�\�/?�����8�މz&�p�΃��_&�y���jm��9?��G��������ix��G�c���Ƿ���l(��0�
��6p�L��a���OC�
��Nǟ+*Z�;<��;���i�%Iq�A�`��V�)�4�4jq_+6#Qb�"�/�3hm>�� h�Rc��e�_�ͮ��<%]=�I�̚�x�]Za�d`�b�۱�ߌ~���Lt"j��h��76b�� 
����Ď,��~T*�d���;�8���<zܒMq��k1��s�a�#���?b��0����%T�I &�zg耉A?�K���R�;3|�����{)��x�����G��|�|��W�6س� �ņ�Oy�?Ο�/^̔_p�lݺU�����gYSr��!������S;-�%��'>���F�{��x��]���+
�V{��s{�'�g��3�G�{m !g�
D��oȽ�w�}VD�y�o���>Aˬ�ʳٔL��I�?/<���u����љ�Ze������p�g�s�>tD���;��"y���70�1�D�0��dCD����G{�������ʬ{1���g�^�k�J��_h�a�Zy���#i�a`":1��׹�|����i���J!!iֿ8��/|�M8NWwG�Ks! s����@ׯ_/o}�[�c��ii�~���Cdh��t�~���¥����h��h=f#h$z��믗[n���	�@0�g��-[�X��Aw�u�) �*,��Ny�ߘ��
`jr�������w�g�nk��{�N�x�K�ʦ�g�E�\f��(�B�6@�|�I+��
������_~����G�h_}�7�Bb�l��h��6RG4ú적~�K^�dFz{�L^ �������ADa��A��W��UV=��������F���
9�A����W_)��21>"#��r�]w�~U H����DL�<!�<|�zc�o��Tڈ�n��K����J�/}�|�ߴn^����jU�h�N���NȘ��o��h���O�3��W�C���GOW����ܿG����㏘G��R(�#����\x��&Pdx���lE��n�8b���Qs����s�\t�����)�V�etx�H�\����4���l-�j�>����ɫo�o���E\(w�q�'&�T���_ϻ�
��G��*��l;�<y�������޹K����h
 Z��H kBҎ��Vc���^'g�`�͓B}�g��^�23�ц!�B7t���o�Ċ��Rq�%�ʚU��V-�qZ�����cCOKg�*ݝ���RW����DE���w��񆛭��ٛ6�k�<��&�|���*�����o5l�!̢�}��_�ݲ՚z䳁<p�vY��G�ذR���ɤ�Z�i�6���P�~\?[S�������ꪫl1��G��6$�B^�}�{���7�2'�3���e�k��h�>�0靣;���Y�- r0������mo3��=��h�CV`�W+E��أ*+�j .�]�G%�	\߈L��O��ب�i����++V�1�Б����,>�:=Q�S^���a1�C���ի�J�^5�s�S�f������J��Svr������ݵk��t�M�;�Z��v[R��&ޯx�+l� ��\>(P=ca���( j��o��x��3�>��C�7�7I#R����W~�W����}��=],����<��òn�2�~���J:$�=-wv����49w�6k�y�g��e+�����/����-�g�
_8K��T0�)�I�VD[ɻ�O�oe�֤�!�0m�ᒱ*Z�����xa1@�Ӫ���+��������ϟ�V�!IZ{�G{���
\둃��;o������9~�������x����qR�<�{X����+�FJDVƋS�C�\iX��{�Tt�=?�W���Vk�T�K�Z��c!!�S^�A넯�42�M���{�|�;�J�h۵�C[?�'����/ ����/[|n����>=�y�<�$vj'|O�A�.l�9��G���>��gL��;�A�S�oذ��;�������-~~X�4�l�֟�0D���dJ��L8ցj��EǏ���	�5�Ԩ���,j�'lT+K��2����ٙ��֟4���0N�0H'�Ux��ĉ=8Y�����q�Xxn"�?2��]w��C�����0��h��;��Qx���ַ�%��ޝ���T�-oy�y�0����]�ش�'��P�̎�!'��Xod�4ʖOѤ�#�$�I�����r#�N�"�(j͞��4Y���ʥK,�a��R�Eƪ�J�%�q�1�ή��d�>�B�%~H�X����������\>򑏘�G�7�����Ѭ�����sj��>�0�[����~������G�O������˭��j{�`ޛ6m�O}�S�؊�M�H���/�5�֫LI����AQ��v�9I�p�(t��XY�_�m۶%b<f�"?�0[×V�/�a���
�y"�Zk׬R/��}�<�G��0�U��/.�JoO��-H�|P?7 �]v��e�>7
���`����"����=��K��?�qz��m��>(H��=컀����{v�o���MX�$y�������ꔳ��,�G��ɤ�,��υf�����6m��v�BG���	
F�X�q��iKu��R���]x�
�,[�R�ղ<��ӪaG�qG��!眳M.�����I\.6r��~`߁���|�8����wZ���ɇ��}�p�c�N�ʎ��q���W�'���ty��"��$V~GRg�d�YB�0�o�1[���,77)����8?�/�ɉ�K�������y�1�_�2�JƻX�J��5*  ��P�����Hދ����-$}��o �?&79�lbC�z2T2��gHzs�}!�
��_��s0��k�:�iP�����y�@��-��y�_����~��,��<4�1j�������?o�j�$+d�X��{:dO'��U���Y��(%K���_n�Q�����]O���s�}��������XИp<������=G^�����1Y�t�\z�UF�p���Y��T���˖�%����bIg���m�<t1$k':>������ :,AI����ÇfsQ�Q��h�gjpsb�#?q�����E�M�E��^@;�/k�B+�\�>ԕ��A�4�����m�=(x�~c�R}�/R��^�7=�`ǿ��կ���ߟ��=_1P]s�5r�7&�W���3���]���j�H��e/7K���&,2�DA��%�B�G�߉ޢ^7�F"�}#ȓ�o�9i��+<���$i$�U�A�1^�\_��WY���0#�a��?���������{����<�B��������0���<�ɟ���gC �y���׿���{��{6Ǆ{�a"$���"S�c�y��j�wȗ�����K�AC�=��/|�K���_�x��s�]�?\,��2��Φ��*��k}�s��z�^t�ҥ���yW��e�^���JZ5m���9�Q���6&������-��A�nX��n m�o��o�{����I�+���bwl�Mr7�W����!�[C52�%����䴾[?e�9���6L�h8f�7+}�
A:��Z���(�sB/D?\}�����/]�tV�����ph�ؘ���&�9ر> ��}�I���JdO?l7�kn��|A�>�LY�r��3O�^j��W�=��q?I]26���
E%9�u���S��ӛx"~��38z�b�	;�[�͈���k��<P��MG���,������gϊ�J?,��`�����C�����dQ���k��mF���d��+L�A��=��a�!��q�Fy׻ޕFrmq� �eq����TM���׾��\W�<e�RД��)�G~L����q�d��F�q�� ZP�<ɚ���7�pú��߿�v��B]f͆�=�Ѓ��s�w���L���zF�����#�=jud�%���~�*&
'Z|X���o!�b���UNE ���R�c����p�v�s-~��
����ϰJ���ߧ�dώ!!�W�ӨI�~��' �q8�^�{���`������8Y�ʕ��?/�m������}�[��l����=��a/���'�}eϵOO�k�ϖ덞�=Syvqs���uB@c�RI`��'�y*1�}0�_��,��y�fS~��{;�{ts�X)[A����g��/�����i�珌o������RR���f\!&Ъ��/+V�2W�O,���a�����zUd������M��0�?�iq�9n�W������l's����xa��%c�rȑ��^�|���� ^�������}sh�֧��I5X�xQ�Q��q�p��S�u����a�ؼ����xp����1i_����5���=�䥳Ё��f��rQXO�+9j9�T*�sCh3:o���뇑�^D�P�B���g�Y*.��(� �<BZ���%�^�'~�i�|�s��yŋ���/s�}��)=ey���>ԓ��~����7��]?>��}$b��Pq5+J�#��a�֭r�X请�[�T�ܷ�LV��l��~y����D��Z�I6?�C�NS���rv�:��\�!~%� ���?����d`�	',V$��.C01���OǌX���f��}�!x�,xp����7[�>� ��O@���͍͌P�� �i����`��%�������7==)��5��7�,T
LB#���~7���$)^V^��ot|,��)@1�D#1�!6�zBPњ�9���0mV���9iı��1{:{���B�����Iٹ{�k�L�/|*&��=P�C��8��g�|�)��1��c68'�p��s�����g���3`�����b`?`��0�9�,{V��y=I���مD�yqo����tp���կ�#����~�~G����)-?�Ž�^޵F�x��\j �B�^1�a�����G��R�Щ�:���N��F����?h�v4n�u�k.�6`E�Ʉ.�ѝ�j����|GN��,X�VD�`#�DՇ?�����w��xӛ����̈́�/�N�`;J�#64��f�Xf��惫⸰��=P��l����D���a�;=\6�e2ˍ�����I,��}D��+�(�yh�IbZ��Vz/��1�ZR�^�C�E��XQ��h>��r��C��,P��J��*(N�p�<��,p*�f��?Wț�ea�8yJ�M����� �`��s�;��|��dqds��� ��1���i��� ���F>�=L�����[z>Jέ��TPիr���A�,�$k0N�Cr�5����ú�0/b����"	,�=91e�	���U���I���p�$q�t�I4�ߍ���X�e�2 ��dŊ���Й78ق���k?��w1|8'��ߩ�����r|�()X��_h�j�Э���q+�D���q|��6�����0�ޜ�W����(`}��l��Ij^+Xb-Y7�0�C\�)���{�� �,H��_=���{�Ռ�3gB��������[�:����\�0�G|v\���p�?>>C�|���S�g7/��J��珠��:#E�%�ߢՇ�b-�o �d2j,�l����&��8�,e�dB��ϲ���{b#h��u��ۨ���?V	�^d}1�0m�� �;Xh�]�X�hcc="��x�ܳ��f�=��C�@�x�Y� a�pQ�R���̑l~q/��(nf��Ru�h?��j�q�)���KH��Й�}V���%��;@ZY�R7��������˾��i��L濓�ϴ9tJ&�vt a������)<�P�<5�����o?gp`�#Wt��Xx�� �\g&��D0֜����3	�3p�����Hl�ÿ*?�M���8����l:cs��17��ʦ�4�e
�,��!�Ű�M|���,�<�߮/�p�=��a�{°�	�<�.����u��3���	�`��&��ǉ\�9|�;�� TuA�Z]zR���w��m�W�@�$��� 7��o�/}�K�w�ð���c0��_���>��ǥ�ǩ=�}�C��
a[`�ִ�o�qӷ��~��k4b���t�7�ik×ʹ�?�8兿�C�0s2�sq������`��ۿ�[��9����p��C�dl�H��!������g{L�F�
lME���j�z�=~�G��>L�'w�3LO���A�������� �+fr�
�f����9�F��D�I�8����6��)0��1<?��G��虑	����d����(L�g}�b�q���sz;�<��6�����Cs���������W���y��<������V$�O�q�8�HY�|O�3 Ny��A}<�`6������b?�O4F3���P���ΰ6B�D�l5���������`��,n��(\�h�}�͖}̤S��1�n�3n<s^�1��;!���Oo��'�s{�c��ii`�u����`}m��Ux'#r�ۢ�+��)�g.|���'�����M�4��h	�0�w��k�w�l��~� 
��
^
@=�io��s`���"�t��|@{�,��Ѭ����_���?}���Ж�-�F�	|�ٺjSP�{|�%ףUT(�ݻ�����B�R=�P����B|�,��9}�d��s�܍ފO[܌��B��z����MFG�J'��Dn�|�x^=(V�2\f?��̦������|�����x�,��I�XC�b~�c6�?9JGR�T+�����������r����>�oQ��lI�l�7\�1L��I~ ���Jȟ�E YR+!�$� �)�1`\0`\�1��]�,ٖUn�w���g��9����;�;��+m��\͜9�-��gW5�?���U+���bZfO�*`A�Ey����.1�l����[)��a�;�l�5�GaY���H(���cQ��p<�-���k��7����Y��{�ޅǰ�����"�{��P�4�y{^[�w�1~�����W� Vڣ�#�}c�+m���?��UuN�W��ZE*e�|Qq�^�-�w��m
c̊;l �����+�u'j����2y��؊S��Y�ąN�*�����8
��Mt?!c��D*d%�ez`�<m��1X� e��8�}[������0Xm��%K�m�p�Z���,��D�sT�����sl�$���.F�<�
���3�56Z��(bKgRzL�Z� ���#�(1p����JX�F�A!Bs��.P�Z�� � ����Fh�ز�N�b�(qL�R�1�B���9f%lR�v����G��9�t�b,��7���x�	���8�}.��sj���ϙ3[Fǆ��zp���A�]~��q��ߢ|�VK��!�дg�A�WD۱�0Y���}�\v��N���Z.)�b	Mݻ
�Ig����uN  �1 @�l��
^�fc!��Z��GX�YL��Iu�����&��N�Q4�U`0��Lm��u,d��dT 2A�q`�)Y�KfNm�V���"��Mgb�:��Η��,��d��r�S��N�	��1��2��Z"���ñ}�5�Ԃ9~�'��ٓ�<�!S�q*
y
��5Pج¦���R����� ����պyO[0�}��h�A�ь� pOj��5HAa�/�OXw���7�Y�
>��,=�9�u.���Y��sf͒׾�5���\���^a���S~6��4I�Ƅ`�g��`yL֟z���Ȭ�3�f������=�ec1\��c����9�Md�6ky���._���b$E��� �a���B�Z�&��D�$�؁��K����d5C
4ݘn��Y'c�8�#0�!5yj�d�8?z�W)Y�O��M�sw��59���ٳba���иy��[�%
�;�.BQg�g��92�����b�3\PL ��X`�cQ� r� b�>�bT���xˠ^-�������G�f"K�L������L�������a��D���&������cl�P"�Nz_�����t����]�O�tQ9!��U���_�����%�8��ݷ�٧䷿�[��t캻���h�)9��c��7��u��k~$/�� �@z��ml�i��C	�z�8y̓/<_�͟-��N����~%[�>+%'�!e+���9&O<&3,ǝx�t��ҎPhG�~lR�?��]�SN9E���_�m�K퉌����$���"2C0	t.BĶ\�ϟ�-�;p΁e4ٽS_�j�\v�eu�t&��Ʉ�&��ǀ fs�A-���.���Q�̟Z�O~z�jRV3�1�
�L�-'ў�`iDs%�0 ��o�a��Dc�p�b}��K���.���C(�X4����C��U���M
e��s�9G�=(ȒZ?^�=p��z��x���S�Źѥ�!a�R8[��>>��kY��f�{B;�3�<ӯ�Tz�rD`3��%q�/c�A��ޤq.4�w���O��|`\<Hm ~���uD�� @;̕+�;!^t��O6��<������(� �z��k�rB����M���;������B��`��� ��YS�  �A�-���\9�%R���}���e��s�;����-�����'w�u�l~�Ey�;߫Z��@�>9�(�t�^{��7����_�z�h�� ��_�<�7�abc�'�	'�0�1�Uc5i=4<S�����8���<�+
�]n�yO��غ	B�q�ʬ���jo��0�?���4��P�h�y�\U�����f�02+�0&`Rt���E{>�#�9s��r��hL���)v�^�����}�m��*��i|=���cM���E;�ItS]�c>)�gŊq۴�������Bj7#��&�׮�S�y��C��82ִ�]?6 ͽO��Z����ZQ{��1f����G�޾��o�J	��P��k�S �,�?z�<��S��9�;��~��<������ʍwEN[�T���=�|y���Um�|L{�6���is���渍}�G�s��;n�#W-��;�ir�ed�_��7�G�B�� �<ޠR��6���>L:�p`� &�@7h�hm���7�u ��6֯����t�n�6H���b�H�9��[_2!0o��Q���vM�ic�Wۀ4�),,tv�����b_./]td�60=Q6�2dtn��|]O���0%�źk+_p>WPE��@ 
��1j���0F��gLJ��͞�-3�5�y�:����S+�A�ҹ���x�Y2ѵ�?�k�
,�Mco�8�vp�úB������WW0�� ���|򓟔[n�E;�q��~a=�=��?%�g��Z(7=	�(�+ȩ�Y����W;
._v�
�#�X#����[;�)W�N{��,ϟ�L��×����twed�K/ʑ+�Ȍޜ̘�U(]��LAd�Z��c�ve��21��܅	�f4�|���Lr��.��b5��XsP+AýMt=�O�m8������l���7HR�M4�z
�����Z��q]��O����y-�O�I��P�4ux�
f��x2Qjy4�q��lf��d��k``� ��x-��6�)�`��ٜf8"�}#�$÷)�d�xv4Ɂ&��r���B�)����^���Q�̙׎!���ϛ�}p�����Mg���|�l�5쫽�?x~�g� pK�.U��������Ö���B�p(��7��`�6�>"�g�d���2w�wÏ�X�hA�����-ȝ��[/\!�3g����e�aK���Ti�3�f�����F��;G%l��-۶=�-HA;F�v�;I���[yL�|�8�S�`�Ϛ�AƑꈺ
�����_�1����Њ��翐����̙77�Y??Lln��I4��t�������y�|��Ǖ�=&���s�E���q`�b����:'s�)�d��]�
�����X��6��f3ڋᩧ���$�;�L��ܺZ@����70(���������3 ��
w�r���)�C!±��êD��fy��6&���঺t�z���?�-/k�P3��q��d����a�ARY�.*úRk���M�m��b>���*��C��MoR�/�� ı  ��s���^{񅗜U��?�(�g���NȎ��q�"�q�Y��ky����.�M�����_|�y�Vp����h�3�Qbb�v�ʦs��Ckԁ��lJ��ɡ��c�5�ӒqǏ�n���Q�ƄM�F�^2w6��d��M�l�9��=a�a<�,��5*���V����O�qܬ`�}um:� �^��8��Ա���}c������cj���6va��Y"w,	0�fy�,X��F�<��gצe����%ƿ'"��®++���I����"�f�q��ʰnЫ�3���|�󟏳�p����ަ�~�/��8]'N��#w!Z6VkN�G6W&���J��`�qp��)�t2���5�6':b<��O��B
d�8�ȫ^v�
��g^�Їv��wҵK���ag��iSK��;�ͬ�X��p饗j�j��@0��{�y�7d�gf�X_��$n4�dL����J܂�%6�f7>c��L���[�i}��\N �1�c5P�l=)sh���8�3�+��
U��-�i�67����%%�k����c��4c�v�9�|>S2Pm����#�wؾ���xnd���_��j��v���������g?��c|i�0#��B����3*�rF{���ު��yi�Q�@]�iY��-�Ҡ����S"kHR�0Г������x���	�_��	�/=��=g�̞��i�nӧ
jrժ6 ��K���\�Grd�5�ό�{�G}��}�k��;�6rva~�+_����7�f�Y�n�6���Zs���u�-cO.�F�d5�fZ0�ϑ<�-@%���Lx�d�Q+4��B�g5|^�~�8s�h�Xo2��˞�ײ��^׎�i(�~3�k����K�}����J���L�eb���e@7yO��ܛ�k��`V���뿎�'�� Ա�Y���cb�
�×.��b5-�l |"B5��I�`����󥧷�E�>�E�B��[+��q���?&o��5_������3ϐ�;v9F}���}��9)�#�fuG�+9YԻ��Ԟ�.+V���-$9Z5R+����P� r�!>����>�1�җ��ھ�ٸ� h�l�7�'%�o�_��%��̈́�ua�sY��M��Y��t3q��2jF�1w���|�y�6Va��V�?��y�ɿ��������
�f�׎5��H��9��[?=�����co�CA`c1��j���]�E��MaGK ��9���{����p�����@	��dՑ�ep�%���B�L�vVB��U�Y9��3���k6�G�@�>�X���$޳�0L��P�����\Z�{��.7��{�L5ǰ��966$4fϤ��v��r��r9�����0�M�6�@N�h,��.�*`��?���p̒a�������,m'�!��Z�e ����2U�:HZ�>�L�j��Ѫ�Ԉ�l�E���&�߼n+���&yV��3
C+x,��cb�Jj�,���P�ot�V,��{.�Z�1Ѽ�m���B���(vC��;3߬0~�ޠAw�&p,���:J��,;���T�Y�R)�M�1�h2�ͻs�e�;�s�tǮRK ���[�QQ�k��:o�WUZ��r��r�mw�+/8_F�Z�d���"�������c
]r�I���^"s�-t����wOp���_���wj��~�� @̶m�����l}���bd���w�/�9��i�$����ؤ�8Y�����h�[ �%��O���ǤO�5b����`�2+k�7Ҿ[y������3��cac��ڠ�T�2�F�9?�ț�[]TlƘe�������v-���������KZ�M�EV,y$s�uI%�{��塇�SO^'��,9��N����]���������b�r�y���k��r1����]�=*]��b�Dn����?�?I~� �'��?��P��c�s_����\�������ŭn�f���9��8�U��� ����=�,���0�9|���*�׮Q낛�n �q�O"^�D���Í�{�I�}���=�s翭��U��H�p�m�)���p{��>R��粩�I����
~N렙�k�u[��<&7�s�T�Ɉ�g�xr�W���Z���fa �?��?W�>g��f�� H��;{��\�J
�9��3�UGɖ�7��� %��L֬^�, �SR9�%��#���?�ŝ5.��s��V��=�oF~��9L��\u��w�Z��	��9G�Ξ[߬nB�ق���u�}/�������?��?>G�=��ƍ��͛b�.d���.Y읤o�L���`l�2�F ɸ,�� �����>P#�ОR��Z�7I�����ͮm�C��7���jF��1�&��~��o����a�k�m��k� �}?p�Dw�2��ـ�����A��
O�������7�M?��gH�[����I'�.���xP�]#x�P��n����:+�?��� ���S|�����^�.`g#0s�q�)�6�}L$.��6l�GyL�=�0���l,�w��ݺP�@��8��?��'�.�={v�;5�v��� �8#i�X�8��QV�>D��`%�ka��}ٲe��|�f=��E]$?���!�ҽ����{?��b;�q��b�
�'2��/bk
(N���=���Nhx��g*�B�z�N@���u�W� S�7C�vI��}� ���u� (��[�@ ��>@j 4���|�Wj��Ƣ @�> �z�ߨ��XP� Y'���
�/Ns���Q0j �vb�:�S�a�#U�C��Z�@�E��x�`�Ŷ��a�Ê��������C? �;aR�g�2�*j�V��R�r�_����ө��N�N���G0�Aq�"Xa���&
�
�Dj*�7Z�����& x!ЋB.��~�a�馛tB�����f! �:�����Ad�eQH�F������Ƈ��Ob�������ܢf�+����˿T�
�u���� �l����3}'����ξ�}o��4SWÈ��aӞ�7���<`pA, �xV2ٌ]@�����t2Ku@+[}���h�$����=����;��&�M[#=��"3�=D��`%��2�M��1����������` ,	��{M�E+�?���� �֮�����[��gS�q�FA:OL�g��|�8�!���Zq���.��-�3+�S6�[ڝe�������XT>@�"�EĎJ6ۢĸ�f��%����{��E~���v��!���p�0����}�s d3�\�f��dVF*^ڗ��BOlex�>�k����PZٞm�g3�OGn'���R� oZ{�z�|��K�4���E��v���_�O�ӊ� ��XLHE��׾��* �o���ЮۅZ?�6����l6������=n�OX��`05||��O�~��/����f��|�+V|L�1`��
�y�@N�{��LZ����'���D�i�	���g�M�����]��N@*=��"�Whְ�̜Z�L>�����҂�}���"J���4PJ�$FK�f~�h��)��ŋ��� �������E�<���5�O�8hNcކ��ֻ�Ѻk��`������ҩП����/�l���m	2��=��f�Y�E�3�#�^����7[�kB�q��>��<]�A��{K=B��/��h�	�+�@�J=��~�z*�׺�ƶRZ�D�02��@<V��oP� 0bҷ�ܡ�$ѯ�ģ�3���(��^s��=C�;�X��e�M|*���y�X���cŇ���@d�X��Np�=�j��e�,�T}+?x>�r����z�����β��J���촞,Vp0E��^)'L��3��� ���ZM��N� �k�]�ijn��1����� ���[�)����U�xR���@�琡ں�d�� (�$Pf�AV�K֊���bƎu��,�m��?����[z��]��]�"~�N��sLg�S�����L��aJ�����[�!�hzІES�g	�,w��ò� N��G�x�z�"��Mz�p��DGc�^K��s�0��շ�yj�48'�o�vl�
ٜf̔��fh�K�k��cJ�RHd��E�ð���;GB'�*��ҹ,L7񚿿�={G+Č�`�Kѽ�:�e�J9�-��0�}G�����/�K�_���71H��t+�Aºd&W���@!�%P���s����O�Ly<{e`�����R3EN[�"#d�5~>�,j�_���ղ��T�h%���󟴁�����5�)*W�:I�5`/GЭ�jݯO���:�m��V�"s�����M�DR����A����YRp�*�����O#�F�;����>;%i����;�̌��B�t���<t�8�T�u�A�,��|���쳲t�ar�y��9�,����NP k
̿
�B�1�ZQ��[u���-U�W���H:�J_��|Ӎ
ّΠ�O&������q½w�*�8>��F�,5��}E�_0[Z�!�M��(`�x�����T�|�[8��dd-�F�t+�L ���5x�*nQ�O�[�,�EJh���i��C	�b$@���ה�����3#n��H��V5���v�I?i^'K��6ɓ�k~x�Ө�ҋ����n0f��i/�]�E�Z��eo�_J��ݲ`�|��;�i@�R-"���4�XK2�Ǚ��;�4�Tg������E(�� ~��3�����	*���䶕���fc�nӹ�̘�#��,�o��Kp;���@�FF��B��2P$0~:P\=�p���&�L L�%���SH4�R?�J�e���GX�z���zu�R�F��z�(�<nw�Z��k�!Ϳ!�}zٰ�1�rMq�1��C�n�u�.����(���}n���wO]���mTQLַc�{Β�YrQ�?�}�i��%g�h�Ϩti�W�� ��,�h��~{�/��Iw���Ԫ���^ɧ�B�He~xǂk���!��.�9&0�"NVkS����g�?W-�� ��T:$�ZY��9uE�
y	�Z��Q�����"�XM�ʽ8U���Gx�LCf=�Ex%fՁ^����
�6k���Z]�&C�X��w�8X�*��4Ѱ��������5p��A�=4|,("+
����n��w�1�Ë��M�����	[���b2�}���G�9F̐l�G��Uefź�5W��xn��3��*B�^Vj�蕙s�h���`���%�<:be�7���9���gܳ�z�%ǐSmdD��i���ԱgYcN<S�FS���	�J�397�9't2��S�b���|�ΠӚc��D���0�FOk���`�׶4���E~�Sr�'�1��؈,�?_+���fb\��B�W����6�ӰKQK�\1�������>�h��[�MY�l(�)��ŗ�RN?�tQ=0J���>�9�u���jr{ٮD�dU��Pۣ���Į5.�ae����$К��������1�*�����o4����vz���hmX�8m>���T��y��s�Nh�Kge�1�.�}%�I&�չ��v	�4CrZߝ���
��sK�{�.'�rRvB�\)�X��!˖.�MO?�kb;4I�4����9�:P�%d�̘�#�'.�Ŝ�3ئ�:5�3β>��3��sϓ�n]A1�
�`~u��ZIL�������}M{���3hJ�ޞ�����sΕ׿�5Z�U.�jZ$�%�"r!k� Z��|��_��6m�tO[���i�j���+9F��c����qV����U  �"�;E��ct%�}���p#�qi�PkN�h��H���tI՜�VH���G�2V��ʘT���v�;�0�B��˘ȔR=5[��-Q�eU�⳺$����L*�Wh�1��~֢� 1,�c�����u2 69gS�|�Q��ýv �Dֿ�72Yy��ީ�������ݏ������w) ��UGʯ�k��m��|��.���D_L{���(f��)��"W��M�Q:��M�T�n���"}�}�`��Ys��Xy��dg�q����ۿ�[\-�I�$����?��?��~���'�&�ැ�>L՛����3L�Q����n仫pH��X�� ���{ѣM�8�B������$,�J�����R�8�;�>K�J-3&Eg%Hۚ��}G_�'�jydB��H�+�Vk("s>@�T�9�WM��+O�������5P��n�U{y�`2c��݊{���P�t��u��l�e�{��J{'��I��� ��Ś�~���mJ�e K�{�ʕ-��P�9�����K��a�ڬ?޳���1�������6Y�z� ]�/tV�}�<�ݼ0.,�#�X��u؍UY���Μ��f�k�<2�n�3��ɾ��x��*K�,��^y�t�s2sV�lټQ~�>y����o��Du��'�g��Qǜ �ן����e�]����s�9��կ�a�� ~�t��o�]���oi�7��Y"֠��h�M�{J��:t�F�J��8���0�i��U�V�-�·��L@�&�]x���>�.�2��Z �4�`Yw���G�1��%���R��ߖi��Z����tYw�M��.ٚ3�L�%�J>�M�`�<S-z&]BG��Y+�b�St"���H�<@� �
{�9�����p��_�=�0 �/��r9�5Z̈ڢMO>��Z��9�:�v�nY�r��~�ٲ�5�,��;Y1�  l��Tb�Ӟ�7#g89�c�`h����Ҷg���[��#����h��Ӣ�����V����}�yH=��3�_ߩ�`,
hӐ�-^"7�|�B�b°@������=��3yV�/j+,m�7�Oj&)��\��(�pZc>�6t5#���K���s�������ˏW&���VI;��7橥*�ʨ� ����^��� ��J�$�6��d۞��m�62(��j{�&�M�&���70��ɸ�M���?�LP��ReS[=K8�N=C������rꩧꞇ���/��b�����=�ZE�ݬ8��ի���O�տ�rܼ�Qyⱇ����+�?,�-c�J�������ΖSן�	
�7>����r��^'t!�)��g�M*|�Y��*U��a��淿��yY�l������^ �<�B�ᑊ�x��r�jY�x�Jx4kA��>K,��[��Yg����������?_@<�І����tM��{*�aG�Qq��|v�P���@Z�5rbld؍u��AT�&��K�?��?A2�j�pM�R�Z��u��b����1�q�5W��ـ!u��+�Ȃ'2���2:��0%�{��G�s[�oߩ�C�c�ȯ�JH�H���%3��;:�&�e1ЦA����*~��R;�1J�C|�d��?^>��O��c���Au����~m����^}�,�x�*�]��2&�f܊*h��wUah���䦛n��K����T�@�`~[p���nA�?'���eK5�6�Ч�yR֟r��.[�̲�8������;�\�J���>���;��|�n:�k�qD��"��w���՗�n��F] X�X�����$�)n{N�l"��tE0�6N �̘׿�m��RM�-��*�28�]
��#�$��|4�ew*]S=� R1��B�3��0��V��!H��ޅ�S=}͇w�x! �P�RtLi�c#���ޤ$���j�I'��4A���?'�4�� �P����:��q~��~}>�ʗu[��x����b�Y1�2|@r���2]tP����	���к�u�E�{� ����/|�ʨ�	H���ʕ��yxý�d�Y�h�����;.М�+����s,�����j�W_�Z=Ǌ+���v��V�m�3�fD�����ӧ����s2:��&bT*U=e�\q&fyX���� }+����I��,6Ӯ]�T@@; ��{��^��0�&:����l�@�|e�@�t&u��$Ԕk1��~���'^>�rԴQN�<&)7���ՃYb��`��s�"��? ���PqO�ӵH��"�Зz`�0���T �� i�C��F.�0�Ɉ��9�8K4ɉ����,�KNͺZ?��.i��F)d� �8X�\�{ҵ���<7����ۥd�&�O���x(rK�.�7���կ~5{Z`���Ν?~�ȥ��m��='�4�n��lA^�a@�c:�1}��}�=���/����W;�0,���k�Z Ӟ�������g�%cVq�3jv��	(9T�l�riDjUg�� �3�j-@*��ɬ��^��T쟋��O�S�����MDs��K����[9t}�"���BA�cHtu��m"�����h���͂^
�ﯦ�W��UV<� 5����%��DA�v����Dh��T�sBp�v�g�����^@���MnR[	�,��-n<�%�y��$��[�&�̶K�G�;��y߼w
�����a,��If�gc}���+�}�ϡн�oTW.��ڵk����C'�w�Ճs ����~��R��}NX��Kh�@JQu5�ᾃ5��R��c��S��i���5sa.1����TN�xs���������� �����G�)Mgh�0����oD���h��Hjm�ק/�M�1�8��h?��f��>7_ǄC���Hۍr�c5���5��w�g.�CuL����!��(����
����gS#��S�o���#_��Pg)�4�S��8rt�(�ã
+h�M�L-�W�g���p5�����M��mj��NQ����Z6+Ǧ�RC��kƽ�p��a�C�>�ǴK6k�����L���%��O��
=���NS����}M� ��e�ݧf���W�������og+I�si�	�2:6,3zg9!��1Z��JM� O{�N���4��]2:R��+��KfΆy��4�R)#]��NW4ҷ��Ȁ/RM��/���1�!��W�*2!R:i���X�h�UW�}�&�d�%�.�OM�����2���̛�)դ�������	c�"恳��+ձ��s"�240���,p� ��F-�� �vL����W��uB�-���5�SH`��J��[T�@� X.元fi�����r26<�n������QAd���t��y�Mx0Ƥ4VԂ!
u��y���� ����|���V��H �:�<���$�BbO	���^�����تZ���x+��o�E�������[������;]W�����E�:�(�\a�޿��䆛n��R�6��4Ȏ];=�������e��Ŏo8K��B�L�o�ҘS��&�/�X�ם�>��%�Ok��j>{B��BӞ����cOl��O<N�֟z����K��]n8!���M�O�����)�y�n9��T���7���>�nL2���ju��
>Z�數Mls�4��B0��dұ�b��N�F�r�i,��1~�؛׮�;7�_�j3��+��(4m�<���������x�1�Z��,��9�|V�n�T��L!�'��Ouų(J(�Jj�D�%��1�����J��r���u�:DQi�Ϟ>|*rxG �>�|��?u���آ��B7���;S�=�x)�������~�2k�B�(��E�9�,��v�ˮ�a9��ӥ��[�d[�<-�7=%��yiFmߠi�bM��0�P�q������Wʖ�7��%-ꁦ72:��9�[4K�=cr����J\,��^zI6m��4�L���ze���C�c �yx�[���e��D�����[<���F͛+����is�7	�-��)t�E널�H�<���x���b���{��k��KP� �Xq�1Y'ra�Z�g'�Tݴ �\r��C.���X4FS��f,�mړw`Uſ����ܠL��-tfKe|��������b
^
�hjd��<�%Ō=ya@!���lJC��'?����}�,=l�<�н���!w��S��d��T�Ȃ�K�R�ʪU���/W�cht@�{�Y����'�i���������=�������'+^�����A��'?���~�+SJer�x���կ�E��Љ�tG�|�4�p�򗿬���1����?�o8G3��

ݲn�:y�Wz�(���3����w�� ��K;w�=�/�n�VՔ���)�zqc��-�1�7`�1e��%U ���6�H�1��z���l�dr�,��F�v�m�]�WoF{�jm�"z[�YhX5�a�k�E���;����d���3&�̝׿��qj7>g2�7��͚��{�Bb�ƍHϟ��.9��u�םr�-�r
�f�UK�\�]
/���s�=�Y�0Y3���Ɇh�QOWs�"���_�d���85nH��{�1NS^�����i�ٴy�j�k�>F�S�1{�cZN#t��-��"w�u�8�%,x��(?\<G}��@�lذA#�H�1V1��%����u�a�d8Y63�L��E����X^1���%$������w&�3�Vא
M=�ˠV���/�Ɯ��%��,��ze�PU������vR)�j�=R^�=�ŷ���yki���K p�iphX7�:��(7]�t&j���U�}�L?��u�?2�Ps��B���ه�d��{�ys溭�-��~��Y}�<�Ѓ�e���e4&�~�z'4f��pEQ�~�Q���~���.�ixƔ�M�;5i�D��	#��������G����n�3w�6MX�t��x���#%�Q��M7��Y���?��?V�����r饗*x2���
�Bї�a����k��ry>�b�����#��p�t��h���6�{ob%��묍�'}�04l�!��2&��(/>����%ya��̎T�U�3�xr���'��3�>�<';�������0S��rJJ��t���������MU*v/�C�&Y�$f ����Q�����5�X �:R������D�R��P�|���hm��×鱳fg�.��pX[8N��s�	���Oʏ�cy��-*l�u�����R=	�06R��z�t}�Qg;M��x≲b�2͂A:&�VKI�1�ǞxLn��V7)��0Y���DÒx�k^����|��؝��я~����.�H���!@��Ru���j�2�L./�<��|��߈����,��b)����3d=�:X5"NۥޞY280"w��^M�����ל�)���$�	��������f����K*�U��x
�?��<�V���w� + Up�A��|Je:�#a��Y6�-�h��m.c���R�h� w��m��;��"�}�yp��0�];�� �p���9��p���(bo�xޝ�~��/�����V�i�3�s���B��]�9�����a�͘5S-X(���v3�]��eǎ��s�7��n�219�D�Ϣ�|`��|,X��H�p�$�7p=Y�f��C�=��(\��	��)bQD��!M�+��^�i�t̠���z6ױ`����Yݕ�\
n����K*'�3��҇�/�dj2�/�
|�.oqQw�s�V�*�=�1�uTS
5S*Pl��gZ-y����>�O~��'��Q�뭷j���ɟ�7����"o�;�Lxf�32tː
�U�V�+�T�`�=�͛6�s��
��JeU��+|a_s~�������QGZ�x�	>$F�ˣ����;�駟�A=)����Ro���(s{Y�?�����%D�V���3�tG�ԑ�j:b����ݡ��s���q4{:=��u*�����4+Q�^��, �U!��u�⎫��X�`�)�RZ���L{��)���x�P-B_��Zw\{a�{\CP$�V�����i�v2-��
�\��tF`3n�v�&.�)�դ[ (��<?�W,�u�r�9x1�����~��T�����;��P�
�7�7
���}H���'u�m�7!]����e�6 ;�v(N���(�5֨�)�u��Ti�R�
��ct���2�[��3|b�KVPE���.0,>�>�я*C�������MM?�zDqd�"��Ͷ��m�����	���)��5�`�&�mj����}��
��_�����>���e�M@���C1W��+��̰V����;0+2D
������(�m�ʒhU�ձ�x�,f����$i2&N�TiV��Q����;�
|�����a��YP������K����BRp�"	�Z�/x��ʑ���u���ǫZ���p�=�oV����2e���#�1�1'��X���7n� �,lD,@��p��#$�+H�0գ��(��[�����ׯ��E0��[�'�֩E�X~c� Ўc�k��{*J�4g���Ƨ��Z�lJV�-?��#d��B������g��WŦ��*�����ݽ*[�`tP|��`��[�S3�ռ���4{@TX�v�=5��A�'�GsX���D� �{��+��)�Uů皏B�.���f#�i���u��g�惻�o<%M�o~���S߱���ޠ��WH�[|�����ˊT����R��~���?92a�����7��.�`7��CVӷ���$Qx�+ΕE��-*�?RG�"��K��G,j͚5��!��$ԠS�:g�&���I'�$K�,��<�ξ]z�]���F�3�=n��A������(�!g����y����{$v����kt�ӕf�(���\�!�P�nӑ���h؉�9�s2���qI~�1d�5TZ)�̮`�O�'h��8���K�����e�Ų�[c��/S&���b��[^����Jf��9\���1�w��}}����x���'1��Jd��] M����?�~Z����&�?iER��4U� ��?��UK%�&�'R}� �糀�����8���?1q��j9��3�x��`m�r����JVp�E�s" ���~V <|��u?P�������O����_��3И��5�-�	9��g���.����C��lAl���0�B,\ &���R��o�y��q�Zf�� ������1ל|��˞�:$���#�v�
���h��&/���od�=���2�aЗ!�HZ�E� ��v�*כ�[�xOt�C�h-
4SɁ��"d��פ�<Y���q�����cQG��e���n�p�?;��x�y�6���.� S�����/L�s&�SS�i�������:9�c�o���8��͟�b !(f���\b}pS��	;aj7�ĭ#Y�x���,�i#��=�8k���� f<@�bQ'��*���@{�>�V��z������RKK��o�
١�B����z\�`��7x4�kLW�:�dĠT��ֱ��!�ݟ|�ɒ&c��;��,$4�k�'
��-Ȅr���wr�;����O� �j�������>�A��7�U2��2a��%5������.K� QK�o!�9�,*�ֱ{O�ERs��x#�_�f��e��߇l��g�}���ek�a܆i�w�駱�t�A�̔?x3  ��IDAT�^b��YٴL2
�yR�d�N:;��e��K�Rq�!2ie��t��h;tY�	�;����e��{A��B�;��ĽMal����g�F��_��EAPW�gQ�2�%��w��V|��hL{�?��'��(%w���b��	Q.U�HWf�T��er��q���S�b���Q۲B�fh�o��-)�*���2��)u�XF=�9��ŜC1�=dD��itD�*�cΧ5O	�^����5�r
!�J���w-ܝ�m����):^�Y��Vp6Ef�6��rkѻ$�Sѻ��lΤ��9�c�y�f���oM*(��1?2,e2)_���	+�5��;\3͘';e1œ~ ���uL���je|FQ��3
N��P-���F�* ����;����K����ɂ�L���+�?,]C��	���e�<V���A)� ��|�7�r|A*���3~�<�fn���$b~���Iiyu�7�@g��bE+q��2����hS�#�[m��G�Ķ����ٱ�������?������}t��� 
�f,)�fY�(�R��|j�A�B�C
̠�3kQF�z.�&��B���|�)�L��g�5{����m=L&?66o\\{FO�2�z���H�g��}���̦Y@6�+LE�ء�Z�z��`�z�S�����l�;d�螱��{�8��Ne��:���;�7v��9IE-3٨[w</P6�b���B9T�#V�/m[.M�ާ=�o��s���DE�:��A#�#��/>L����64]wf]��m?�mMlLl�v&�mۙ�v&�m��}�u��9g��]�]]���[g�֨ ���p�Z�+(i���Tߖȥ G�M�qdM��2�0'��^:x7-��R�af$eS�[���"*D_٢U����	�&uj9ad-Gv%N(BJ�J����
�ǎ��B�wh[��zZ'.u	3��c$��6:qd�l��&�%�#^��V�z��˚93�ٷ���g��Sq|ܥ	���ʦ�&�8Iz-/@<2��TG���<�߬[��X�j�jZ��U�������q~y�J4C��h��"]�j����R{rU�R��4ǣ����T��9��w�Ļ��<q�;�F^���.������LT�"� =����<4ƙ��+�����"�+1�>��T��$-�*��y�D5Vr�{�l�:�r�Ԋ±�Ey&�����1��d� u���b>�ѐ�N/�7AaU��R��o�tY1�7㻇X���pNcf�Ov>6��þ�p��wH�\��lI�`��I4�+�=�J��!p���s��ɰ�F��X8E�8�SԞ0o3Ĳ;(�w$�J�0�'�%v���
������ 9�:Lf�Wew���c)����p�"Ϟ�Ê����Xag�5&A�H�� !O=,��{�s�Лπ��.�ga#6�J�	���������-�%qH>Z���ϗ0_rP���R��٣�!��H�֛�P�E���7>�ic�����v��:w�:�I$W�kj�o�*w�[vq{��ͼDM(��ʗy(�S�}.�AO�?�p�����i2 X��MB`<���P9:�1o�}0h����6wp �4�\t]Q��@
&uUS:F��f�fD�*��y��Q�y�kSnq_�W$p�^�����Q��R����^�_�<q_�e�}�B	���N�o[3��!#b��V��.�e���	�Ȋ����~��e.�a$�j�\k�����l:�a�K�8���d�X��y��e���s���	$X��D����Y��S���p�?��B�i�)��F���Y�*
P`:RQh���e>��!�mN8�Ev��q��B6�~#����3�-F��������2�������ҟ� �R��U^��~�+�^?p�������濑B�����ݗ��o˂Y�Ws.a�J�b�Q�hT��'�]��M36�U��4C�'G���{wj��r��F���!`u����y��)U���>�a;����f#���UԚ�H6�뎛*S%�;ڼ<��3�Y<K�6��������C򬷟���d�=w͌�c����b��e��q�(_��1'@'>+�>�]�@���m2�ΜY���c*�x�z��T�S嘎���Me���Od��3ǔ���˭:h�l��1O�k%��S�:��쬧��SZ�ݾ�]?����S�ܽ�E�/�	�\4�M1��6_y���d�j���Ue1���ѐ��Z���,�j+b�4W��d�aɞ���D�����qAL\K��_@�q���s��Zn02��k�4�\�k��<6̵���[+&�$� �>���k�������� wf�:�V��>\�e���x�����*�;�M����F��g��K��;Lyk�����Fe+� 5iQ��.����4�������/1����Yj�4n*�����u*�֐��P�ɿ����w{�����ϒiF�7?=�h��.�bW:��Z��.�� ��U���ˬ1�x����Y���Ԣ
�W�ߤzB=Y�B�^_{��9|vڤ���%LuyU�e �-r��Jڷ���n����(�8��rk6��q�Aec�\�L���o�*��DP�m&O{y۹�o����8�3���Bi�H�~��P9�������/�*����3�%�#nR��ViӞ^0g�>D��,e�T�}�:�9�i,&y2��^�8x�d���4U�pQ�0��8a}�K��``������F[�2c�K�QW�n?���9�>�~?��nkw��-��������}_��}�8>�i���J�� +��L�=c
�+�X �kdw�4-�
ʘ��9I�b?F&�s��ל��本�">�IoL检�*Q�[|�ɖ����c����8�&,G��d�}wJ5
	;�#���q��t�� ��{�P��w�-a澜U�� ��@	���?z�˸KN�|�}���͜VK_�Q���?����ZE��~��}�6[���f�f��ߟ��U��0Wv���c��Ev��Q�	�YH�"�W&�W�B�xc�����RkV5�-��x���������z͊9[w�<����e�|Pi���R�<��q*�,p��*6�n������&��R��q�
�v�s�z�q��=�Uv��u��\�'�������i�H@7���I����ӱR�V�֋���q�$�+�Sw98H�t"�y���ݳ�|�@�ٴ�p�+Ŗ���P���u�m������Xzl���Jp�� ��B�m���=%����:��"������&k,4�}c��I KW���Y1�dx�O�ϓ��zM�>�zUn�Hv��/x�6�XE��S9�	O,�����PP"��i���(BZH�]l�n�"�Pnr0�i���b�o��$�Ѡ�j�Q���T��.��Ѵm�~�1>E��浱se�2^��$��w1��P�h2�Dt�oh6y��:ltL�3}P��<2����t�	�/��N�(��#x�bL�����Q��?0RI~U��?&[g�3A�� �M_F�I}7F���}a�A[m�/���ؠ�p��o�qD6-"'�_��t�_O�ze��sT�妅�t[ބ���؂v��~`��Pq�)�)��&�鄲�~�2-5ڐ�# ߫�D[��QH0�P��e~�Vy�I��C-�L��Lnk�6�a��s�7��}օX3o���b>UY�3}ف�u��ߟ�V� ްU{���@w���C�t��t^��w�*�gH���Y{iǑ0�\��~X��6�:��!�_6[�Օ3<'lߌ��>���'X�&Yy�4xOʕ�5�M�iDc���`���k�`�0qA	�7 ����I0@��w@@���'3��: �D��q6Ap��uX��R,�7qş� �N�����9{	#v$)�8���Z*��s� �������=�[�9�[yK/]���ZI����.D�܂K6�M3��,��r��G�X@lv]��.˹]f�S��T��,E�pQxོ͕K�m�'o�;7��\�1!2z_w�lN��������� ��&����v[�a����Ƀ��
�d��-J�����,�vUP�?�Av'���/-S0d�����l�2K�A�ړ���u�N�咕���N(����j]���O+"٧6�<�O�7��$ޝ���L���,^!=60��E�9��}���agM��%�O�4���b�ˁ�^b�H�{
P눻�#����v>iX3��#W�^3�_I��r���I�6�lc�����p��n�2��v�����4(i�n�d�N�ˢ�3ރ��+���Ӏ��řp.p���c3�]�b��]�5\'0���ۦ3�C.CS�k�[Ҋ(>{O�&1t�/��ȹ��f�{5'���Ϛ&h&���o�^[,.g�t4���?�cbm�P�%����X��'��ۧ�)z��
��7^��?�{�S?w�)LК�;Q:�3�z:,�13،J�toI�J���{7&1Y?���=�����%1�ޡ���V�p��Vè��M@����8��_����A�V�F)�ĸ�ު^�WՑ���*�.ܙ��h��c��|���DlJ�S}Π��ӊ����?m��,���T�&�%����������{�N�m���#_@Gc�ΙA%x�����6ɸ2���
�e�;���,��u�2庫���������~a�/x�IMyHvVb9�6�^��̨(\��O|�*���t'�l��U���=Y��?��P8g����^i?�o�Xy��3�"aZƟ;XGT-Z}����wy�f�o�侓-��Mq��lL0�R6d	�_�V��1$���i�c�OB�0a��� @b���2 ���i~*1���/�/I�M{�����O��_�y<?�xJ-DP�����qrb�G�ǂ�������:0��D6�:($�#���%X=�il	q��%���}U=�MG*/�~?�.�WQ���^w=��,��$*(?���.�����!Dq�*��NI�<��]�ǥ�T�8�7,F�i�����\�W��x^���+7{&����<�`��;@#��Ϯ�,h�/�s���K@��e���I�6U]E-�pj��a�58^$[-�3��.��e�$�������!ѫ�l�hO��91[=պ���\l�&@�u�2� %?�DX�s���bYow�����H��i��l�">V����B
�+0�[�GAKI8	�m�[�@�Q�̈́�X:Z�X#�O|B�@X�^���xwh��!M���E�q�QAsJo�e/гInv�{�������a�(Wi�5�>ig����}M:��=��b���W>�����Є�De����+TǇ�	t>;6�y��l9�F��v�6�������W$J^7K�W���`!r�Q}��%��ƶA�� �q[���� �A���M)�]�j�v���C�ڂ����ې�oS���bg7���C��|�خJ��}�h�=u?�.�E����Sr��T�ݸ*{�ݿ�%<:j�ܹ�o1i�y~5�Uq�d�D��kf���_�rAc�����śᅟT���I�}�a&|0e����?�6WN�t_Flr����1�y���?��(��f6�����7�[l�Gr#
��I+7� �Vk2~����L)��z�EG���x��W�Ӡ�~l ?�-ؕ(����Η����2"�2���ԩ��a�������(�Q�ffe�A1,�f��yj�a���5F�j=���^�ŃS�_����{|��ҎOj/ ���=�p�6�4ͫ�B�+ͬ�`��[q�MR�Z���S��gt}u�|X��2šT�W���#>� I�C�v�-�r��l'O��__q6V���N����Gw��1��x�����y���pP�Ӝ�鞐��ogiVģ�A`ZڻJ7�8��z^���H`�L74|������6E�P���GJ>DJ/\~6�]M|]`2P���q8T���lF}>�g�����6ZlFe��M�2�´�뿁�g��c�����Tڽ�z^�������s,�����|2��/
 >0�����mp��D��V���#4������ G��4�	�iC��Ԓ��tR�L������P�"�
S���ڷ�ڕ�&��<'�����{�c���t��ð.���Y2C��+r%̇�f�<�0/c����k����և���� E/-F&Pɫ�{:G�ifm�T]/����$_#��s�lBi�[��^���R�Eb$ZiF�(�#�TD�4x��F*�$�����p}��R��k�X���n��E�Gs�w҆�<���=��͚��;����e}Z���#̾�!4���)���	p<�v�0K&��\�M"G]Z���gf��?����%���7`h��.�P����m�ҵ�}v~���B�4�����Wg5���g��|6<�f_�=�i�;Ё�t`W8`}�� ����Y�۝���^f xsL�=��Y:��W�/�2햌nr�r�w���R�A�[���T�b6N�m�X>�6�.}|q�Εf��MPl�O�+�Y���R�oQ�l�U�.�H�����!8�'Fͼ"�EC����)@K֓��lY���q��H���;�^�r?+��/<տ	>Oěb ���i`�n @����`�!X�~�AFepB�04<7H���Fh�ܼ�iC���$�o��0*B`��oScU�<�K�*��8�B��Gi��'{�"��ί�+&B���V�`�j�����& Ͻi��*+�|���4e9��4a|�����������93D��;s�*-9Uܳ���$P�O�����*ίv���!��?V-:Dq�y�0�O�G�<@_>�nyo�X��D`;\L�9����xQۂ}�;T~��V@�(��4�ܰk�>��T)��1��?8kMi��Z8?A����y�D�!8�M푕�4����s�2��29�3L{>��q��3}z����8�-��L�Y=��@>�d�Eq=�BZA\\�s�;2�Zqbc�\�N�^ՃC�.�r�X��&\��ό��Q��@Eg�����DW���+!$1��P�O��9��ʟ���	����q7yi�u"���53Сz�����bs��U�:�sb,���˘\��W����!�{?5��c���Sc��y�:[>��4��Jg)�l��
�M�r���(�����&��b�@2�33�͠Q�Y���!��U����e/�\3@z[�5��4�+��MUnw/>��J�\IY�׃��z6E9<�F}ŭ���2K
��?
_��������#�lfE� #�k�^�7�&u�-�A�{5�{�ߞ�**��rI�$;=;�V�,��Z� F��/Pd@��<��6T����w��p� ���=���)�h�����'�3ٴNr�d��8=}�����Ue����?����k��t������G~�@�`;}a��){พ2ki.�R|[-,z�0�V���ex��/�2{��.D`�6��t�G�.��?ו����&$$�(2���M��l���O��2%<y~�,�s�I�i��;:d쫮C���[(�O9��KW����@�Ԛ�ݫy3nd\`��@�!V��>�XT~p�uá}sam���!*��F�� �B��2.���l��,��ȋ ��§[�7�~�YD���yj��Xn��Q��Z��ct
U׈��.�^S�g?/E����}%�	F��z������z�:���8�A7�Wg��2ݗ�E������d1z���T��(e4�#���\��a��쬧�<�~�Rٞ0e;6>�cO�8	����f ��:�y5X�R9��[ۜ?�%P�}�/�ҋ�	�Ve��]�t��!Xգ�[c�����k���!�th��c\m��	�EE�f��v��2G�R���5�1�π�vR
KJV�&2115K�T]Ϭ#I�������O��PRel1�&�On��N@c�ZcI�)���J�6��e���)��l��"�H�T�Q�V6�`ɼ&����A#��e6�!���<����Q�&;g��X��X�P*�+��˳"FOX�+��b�!L���Րd����(������p�G�.3�Uƌ�0T#f�/v�9�թ��0��|�����^+
���ud�]�,�)z�BOG���^��%y�=��'����i��u߅�*�:���1�i�ŝ�J�Tń����6 D���@�Y����&����+��(������� ����3�������L��DO�%+�½d�W�}R3;c�=2V�|��[���
�c�.�yf�B�BK-�X�А�s��s�+����MF��P����!NK�B������x�T�aӠ�Zbsݞ��:��e�%�;4�p_�v�0��ÍH�X�U���{�pa�jbi#_��	RԩybN����N�H�߼�y���"2��V���ui_�����k�X�]j8��w������F��~j{і����5��Ԅylze�S�{�P�P�9q��x�ۦ��Ɉ��ᶉ�ځhP����8\���j3g�K�c.G��h3�*W�a-W�&˦��/a-�Ȃqm~��CBZ��f�k�⦩E�5�A��10��h��&��!S��q|���t:5Lh�<8���P!�vxӻ��U]{�y�7����ЩyI��k+�&u��o�f݀��,���41�����;U����˴)9�q�1g���?��R��8a1C]����^?a�˶�� 6����WMDA؂�֟Ɲ�-�E"�W������������Ǿ�8�:��=���i�o���������|ʩ��'��,�vz�`s�(�J|lG)��џ�|u\�S��2����l������r���#.[�m9�<��%&(f���]�"#<R��o��X��1�ϥ8}�_'Mf�7��G�M�ƌ��j����*s�PR"3��	r��S��m���X����7��+���3SbV�	{ ��+
�fN��v���/�����/ΐ��Wl����SOP��_��|�)�ف���+t ��'m;�W����Ԕ'[Z���ο��h������)g�,Or�}}����~�]D?��+�fu�'���R������t���lን���< P��k"��i����jND�����$8oњ��ǐ��a��{r���r=�r�!��N���� ��Z��=�'�	��7À�x��vs&u,�Ѓ@��w����VʀS���N�)���V�h��d�C"�ĭ���m����y�7�@�N;��G����(�P�*Ćh�L��6�������;$����ʢ$�;�K�2g~�D�\�qUu�p|�*Q�]�5��8�	D����o�Yf?=gD_S�o�	΋ꮇؘ���O3&2Vi(��:+u$3��&�ځi������h���"vA'�}~,���sݏ�3�!��0����l���Eٌ����]&�9Xq�$f�]���h9`rM3�1��l6Ĉ� Pʔy����(PW[ n����u���m:6;f�q���7�0 ���B���F#�e_L#-����414.�sZ���0֙�`������VWd����kc��N�vӜ�x���
���z{Ðn�R�ya�qE%��r��q�}�,���L�j�"W<(�U��~�]�giդ4*�Wo<k�~��E+NР�g�>b�f,O������c� <�X���� į[�ѭ���1#~	ڞC��x&����{�M��	
&�d�|%�@'���^̞���"�!�|5 �	����V��y�z<�(kN�jj��p��>��`\ g�r��%�A ���y+nM�F���|.���{�I�L�-S�l�%z2a�d�f<��ǋ�<�QxY�	�%�'dn�K�-�P����֏j3�q�g�2ܿ��Y���1ط�Ƈ����#��ʻ���C:f�+ڶ�5+��C�H�ge��������}Vai���j�@ݤ�|Aw�q��K��Ҝ54&�ɣ�����)N5������{����4m�g��(`X�~r�H�H�\�����S��+P�4��ЉhM@��N�*&��o`��L�YB�����b���M5���"��׶�Ҝ��":�� u�'��[U`�_^��>_f�U���\�,V��������}Yu[
�g����a[?7��n������n�r#������F��ϣٮ[D-�O4�'j����9�^�E�O���:mwHeKB:�J�']#��e�	-yGK���I���yg�dm�9z�K'�x�����,<�t����1G�؆OE����2�:�Tj"99bDE�w������m�f��m˳���_m��1�1��Z���G<�@{kK�
.Ԩ�Eۼw�d�ctɾ��%pƃ�b�~Y�WTk��-c��
ED󰘆ou�2��]צ#*�QVK0����b-��*I1Ê	�r�+�i��1M�
9rU�hL8;�;٫�����c�^��ȴ��������a���(�}�FEiAE��h�3k�����faF���M7��Y����|�,B���)>�^�E�sU0�1_�	qrݴC�!�o��Z�2�%GRs]5/�X�]F�&>�����AX�M���g��P����[��:?3YLt���:vH{��R �C�b=%VQ��sa�^X�<U!��a�o�c������9��3��6w8v�"�Q(�\�B*�V6�\y:�ߗ�#M�o��4�>���ګ> �څf��� �����k��^����MW���p�N߸��n����A��Z#����8���ԨbFFn��mR�y�W�ǵGA� �}`���N�q�R*���L'5U,�ċW�L�ZiM��wծ#N�|���f��*�j8���ru���g�����ɚ��T>n�\��;u����q	��Ǆ[���_0FZm0��K���	���:EH�Y�G@�O����]=_���T���m�r2Z(zz�(E����>��ִ�o쨈�U�*���B ��[�lk��r4�-?��t��8�o��+'z�C_<�3�� ~@t����eveP��Ui؊#�;��B몀�^�-��Y7�:~<_G�E�*+�j4�G������s�~}r5�A� sq��z�������[��I�c�!�vhJ�����R�B�4��@G�c"�f.l�����jUbA��ݱM�����hz��ǧz�t�E��醧�N8p�!���ud��s4*�}"��b�Y<�6�S��`�����$C�(�JV�#�QD��e�TG=���W}P��tڼ�����&q���u��>�&��ڞ��dY+�|�)����&�D�_�4�L�Ԇ��9{��k��'D�	+ۼ��4����0�~��hd�u���g�{����xD�w���`j���0�(��~�޴y�Cˡ�ތ�#�w8B��!q�>X,ލ�Vz��������O�V�P���v����5�x�ٔo�rY ��&%d��X�qm/4#�PԤ[�����������K�~�V���a ��%��f��f�l�y���g��Σ��TR�gE�.�m��-�)���M�u�w��Ix�+�*��l�+�iSD>{=f�X�
/f���V����#���Ql�>���6��j0��5h��E�~��a�����z�W�����M�f{ݪ�JL�tqp+wK��]��觰�:m����2p�H1�q!s�3!9�����u�y�k�/��XZ,s_���|��Jʋ�k]5!�8�`�e�Ì����b:��~'��Nu����ʍ�ڻ�(D�
�8�x��܏�G����U��J�Fa	4j�i�`����1�L�f�P�Z�YOxĘ�B'�?���,��S�D2HR-�_���0�����a�F����jn;�r��~ʊ�Y?�Pފ��#�J�&����pe�� I8oo4MkRp�;�4��,��S���ͪ���l�����Ѭ\ ���Tc�H̦9+�R'շ7�����8���Ź��A����A�2(���F�\�;��!�4��ܯ�܋q�O�%VR�i&��!1D���~+��z�9���i���j9��_����V��0K�<�3[�9[����� L0���q�r(ڷ�m<t�φ5�=�!P��(gN�^*F����d�GN6ĺ演�Q����w˧�ޏ�j�Ӷ�Q���4�ph�L ��	��w��1����ݝ��"��.Y���$UL�R����O6߸@�=����X�˖F��@���R�!u��v�+� ��x2���(���g�͸ �qZ��P��8�	ru���-�#���~�#>��3�jC&2�@ӟGv�C��lV�w>����5UM,��+�4�M�`�h��R���4���..�I0f�?�,nT�ϖ�>4�[�<x?��}G�%U���0�D��0=馒����Y�4��t�lF������ ��k2R�Ԥ�^����GV�~���O�'�Ŗȁ{`������?=4�RzخAI����\ZCEj�ϔKϡ���_�sUX�$=�]�>;nfQoP���({��܀�l�H��՛�w���o�&��_�Aq�[�н�Iݟ��kxG����wi����F�B��KIh�o�S�Fo�����q�7xz[r�{k�˻N���@wN˂�+{q���Oui&��*ٸt#�LpŬ/���L�5���W��xبN;�W�n�'��*̗���֞�����1�*�ZnUt�h�ZӰ/ǳ
��/R� ������P$Ɋ���d�f��,K��Hj��Ll�rQp��:69������gi�c/̷�Z��K4*S�uוp	�땮qY�}kϛ���:���dD	l@g���#��E�fq��Tύq�s����KU'(���Q$��t�zws�"oh׉��F(V�MC��x��j����+Ȗ���5�j����?s����hu�,�0���=��\}=��d�
�c)>�&�����d�칤�]mҐxc^��V/tE��}t���aT�gn��~���kͪ��`����X����h��|��QGb�{9����E���cE�Z=�U�����Ø�C�C�e���K���k�0"6�d�}hʱ�}��5u��TǕ��G��\��A��K]��=��h�]�l�E�[_1+��Re�Z�ݢ�]ã�m=�]�,���
��]|l�coyiJl��	ǖ�1�VN+E����;�7$��٣#�&��`J�!bh�^���`�����IlW�0���W�3�ƺ/��q�b햢��ũ:<�MS�I��os���L����qFv��~���aDmlp:�Sۊ�pU�0���U���W�NC�d�t>I,�ě�����j��usi�O3a�1�j��gc�Z�Y�y�9c�U��mh�!�7 R�e��v��W*��<���滻J��\FrR���b/U�����*d]g��M�B(�K���L������s��'�(�A��&��=�����G��_ys���S��rW5�]+���e�J>��vI��.��MJ͒JM���F*R���[���f��+d,|Qee�B/��=kx�]���`Ѫ���9��uCX߅��k1���-y~�%k}�=�@�x�!p9�g��=��́���!��`�����'瓮�_�x^�o��@��'ұ;�u�D�oxS�rY�k�0%�g�^��>�h��=�#.U��_ay4�}��R��F?�J���}��rq�D3�BN�:���[��$���o�E�����&��d ���s�z.�7,"��������Ie�9��J2�fqLR��ņ�&�:�E��{���3ב�*���ĭJC/]��fd;��,J���\���
�5����{O�H�%>�O5���ҁA+�m�mB�8$�4�e�*}�j+�)����{��s����g�y���7��r=�z�S���pl�rϭy�z�#�׻F���[/�/f���R��m9[s-&�1��/R�%��l9�D���%
h��e۰#�u�kB��t�reM}[x5)q� '���sGӵo��R�n�|��"��)�{��;$Ӷq�m�c�Y_A���F������k��v���O�nxLg�m����"�3�*1�Z a:���I{�L��Y���kX�5���-�b	�	܃44�R�<R�׻�4؞�G_������#��͉�a�;̘���l4�ݩs$��kͮɾ�o\��� KR����v��3T8D�m꫏�Akc��TE�n�u�}�@Y?��}�� y��Z�4��c�)MG�ї:���=\�c��J��eV�� Q�	r�뢞��UʥOs��꿼���.Еo���z����t&���9/G!GJE���$�cfb�t㻗��b�(���Nɧ{�L�²��$ط2\{��	X���<�8��C��1 ����J Q�L7u�_�n�3 d���C���ݻ6�:��:���0����<�K�x9��7����w�jZTn��&�9踰a��0����ǋ�T1�����@|���8ːy�[M�Y����g:V8ݿ�f��F��[��r[�G���p��軨�y��˷����QP�ˆ���mu�3&Bf���o��d���0\A�΄V�@Ƨ�����Ӓ̋>Hg(h���Xg2�ix���}DO�4m�x%�̌H�����]-�?�Idր:NPTP�\����5�l��ѠC�YC�?:����~ޠ����u��y�y�8�$�;�+D�8����c�a�(I�h�c�;��r(Gcs@�ĵ]�+���%�`�'�>�#��4ٮ��G=��h�W��Ψ���~�~kW$	�q��x��.��� �m
Q;�V4}��,Ű�;��j�*�*��K�I�����������?�X<s��(�v����ʻ�sBA|���1��oY��}�'m۷2��f�V7�43��X�m������R��y�{�tbh>�CG/DvP�C�M#��O�at��dy�N<�ȋ� "}���L}�0�)f�� ),��0:��6C�Ҵ�N�!i����Q���d-�ؒ��x&~..]R-��/��e.����b�[�E&+�{;۾s?	I7���#P�ߡp��'�{��;�~,`x������6&Vpg�F�����\Ы|f��3W��؀��n�il��Aư��b� �j���f��k��92F��.v���ya�#I�g��m��_�*�����P�ߕ��a�^<�89"�A~*��J_��bf�Qҧ)[�i�V�+3*�z��*O���2�r��y��m�i�<,��%�྿7�Po�`�1(��O-S/�X��v{�M�]sC�zw5���Yt+7*Hb�㾤2�À�O~ZЃ����m�>%/�ZyZTw)k������K������j6��~�~>��b�@'��35��hGAB���ß�r�k� ����N�h_D�~m�g�"�$\��\�/�A�I=���\Da+���������Z�W��%�ʕ^:�I9����ȷ3eE��6�lRҹH�@16�L$�P��Gn�?�W���kh2A�^�g��$x^7!�&�������� B�LjA<��"R{^y�<��<N�U2�z�Ê����ɚ[���V�~:+��}|w�1���_ݻlߜ�XY�B�#A�,�1���'?�I4�S֝��3#���}�ヶ��k��ֹ�E! �T��?Th�'�/b�]�����R�*Vx��T��uXB0o~ ¦q�"5M�ɫ��os������%�(�Y����FU�����/��y�r��DѢ�J~ �t�{=�^��$�	��#�_�� ��E�ơ7����ҽ��#�EFn�ɸ	z:RU�oxx��X�?�06�oZ,4p��XY��~���	
�Ӈy9�%HkĄϑk�O���79� ������eK	��!Reo��a�'[l�]"��%��$�(�)A:�%����9qRl�{l^,��<r�-_v%�R3�J��2�╌'U�Oבb[�G���8�
���7+�fء68�ɅĠ#)�B��2L�6e�R��}�>Q��"�V��g1G�3I0f߶�qݱ�Cς�c�7VOS���ŬM����cy��Y����!B���ɀ�1�1�����v�����ro�Tۧ�����\�4�Ut���֣�g?��?�����\#�>�9� {���K?����s�A�����`�r��u��� h8U���)n�Y�N����R�]h�*��*�L�+�m}5���+�_��%��*u���E��9F���y��a����L.z�Yu|2fͮ�A��&D4�Z#�)�<"��䌦����'�&�A��xX����oӑ���I�FB���������5��|��0zw	t��7�N�m�{�仐Z0Z���h_����;��w��`�G��T8�O��������rZ����c"i!X�����Du~�he|�T��d�E�3\������eۏ�K⫻i�g_���ޅ|�c���mqY���Ѵ�>�*8�qX�ȠZ�f�|*Ԁ����O1��Э��O&��qᅬ!�^f8 �b���]����00�xՈz&S�HmXkU��~���w0>%qP�U8Q�.��[�*<ބN�v�Y0���xdg�����4��#L�kh��.�4����#^=Q��6�
9 ��o��L,�ߙ	k[ͳ�Z���l�CIK��]��=�zN�V3L��<# �6����/}!�(�QN�R�Gj�4ǟ��n@��w2��
�,cջM� �cRxB�ݫ�,R#)��W�m�����}bu��s��(V���?	r̴%�=�1�n�&6K�_��ˆ�=�6��Q� ��0�����%XĒ`0!W�b����[��G�Ə��=�5=&��
���pL��}��a/���!�b���H���/(�('�,d<��hϏ8�0�b�2�ڶ&dݧޛ�s@T�H+�$,t��2K��G�X�^EMcFv��d&2ۂ�eYM�8ZI7=In�D���7,�'\KXŐ��qa�6�^���V���.s�Z���t˜S}�����@��#�b ߖ���it?�ca�cp�_�D��"Q0�Ӏ�*�DE˴���qA g��@��a��Z��Jd`�d�X
����bP�W�4�����2�!H������c(��hS��+Z3q�U����� w@��n����\OY�LADٔ[��fQ �L�Q���OU�2->�ӅvvW����4�T�X�Ey�۵�F�  �Z�v��V^���Y{����Wsº�����
��xd~CP����_��o��%�y�J��E���s��t�Iv�'z͍���f7����,A,��/���Dd(�AA��Z߂~�<&�D�%5��<��|&a�����`��]۠�2޲�y�t~j<�9~��G�?��!�9�Aa����@(�L	�~���g��:7L�/�����u
<
R���
$x3���y��Vt22���KVy}j���-[��p�p�1�Ⱥ�{X��֮;2��<�kj�nU��=�=ϩ]�O�m`�f[�n�]#��Eg��������wXc*�����!������#E���	���z�B�&�C`-!gT<R1 ��5��>���;�$�9x�+^a�������L�=�8�ą�llv���\�M��#�o��j]�!2�r��R�����G�M��N�`3#��f��M���|��ށ怍MYo}�rJ(�E� �α��T3L8��K_�R�`�6�5���aY�z���\*[<o5ptʔ�n8,�V<�%���_�<��4��7�:�vf����>�-�3r� �+{��m��͙�O���3[�G�-�G��jj���P���d{hƼ�E�r�adF8�9�}���۷��-74y_���}�Z�t{_Z�u�Mo�2	��]`�Lf���X��h�Vv�5��cc��z��|�� Z���B�O1AM��!�������P��[�/n��-�#��=�	N�t��!�ʱXt�1���!!�b�ϳ��*��k-Oc�m@$��!$��eW �to���ޏv��ɺs��/��pZoI�4�lr|4}w�W����񬍏��/����DBXR��{3�\����,��莴Ӈ�w�Y}")��	� ���Ζ'��{��~�j�P'��C��/��,Yk|���kr���it$��);�3=�り��[�¿��7��u:N��{���`/������$O��g�����=��cNGcA���:�l��5���Kq��|��ڱ���Vڐ�)�zc��}��!��s
�}AG��-��`�}�L���y>b��#.�����0"�0B.������9��KC��]��{P��W�rn?�!��7�e�gX'S�j�6h͵����*�{+c�����~���dm*��]����G��~��Ie̜Y���=z\���G��O"�/��iC1�\��U�����{p�~Z�>zZ�s戮�?fc�۝�99Ѱ�;��W������^ ���[y�,S�L�{���66���$ͫ��t/ɣL
��(�t\#��N^��K�FQ��=���	.���l'	��K;(6����l�F�;�jW�ȚfRV�&�~����g0�>�\;㌳|--_���~�/�Z��[=�����z�pݢ���Kie������<+=��/�'�x��=i�֘�x��~���i�G���k��u{�K/�3�8�'��LJ0^%6q�#�8>�h��y��z �\&kQ��9F���0�s�(x/�|��f�tfs�����+�'E�8�<		љD�0d��#�,�ى���Dƙ���	2}�����"h.�c]����'�*g�9����SXO\O�qRP�!�JO��ݺ�lw$���k֬����:A�48ɡL�v�u_K�`�v��Q+�j�Z�CIy�%,�q�fV�U�
��u�s��DY!���R�>b~���M�/��j�aOm|����$�������Z��{vϝ��ӛ��W��5�`�,�+���6=����;�\�4�^�[�'ּ"�g�y��Y��v��e�n�d�c�����Aa��Z���i�sɲ۽{�v<7f�z�o��N;ͅ<�:mv�8)��đ�O�=c��G}����SP��^h��bzc��a(��"E6&�D�+:^��oi^��
�J(K��<���{��X4�!�ň��D4}�<���P�U����,&������,�邔�o��	�$^5���=��g���V�В�[�K�,K�g��O�ã�+	҉�,ڪ������d�����7����[*��wK�Sʼ�bm{�(��L#sK�Z#����#���_�`4�~ޒ����lI�'á���NL5l|l�x����/��b�y�a�=>əg���9`�����F=��Sltt��4��v;��c�ϱIP?bc��aU|a�	�vW���^���y�l�&y�{��]�轉r �o��o�k�q%��_~���D)�S�_����z�������S �K�ySB�	�L�
D^�ޏ�:#�^�}��)&��K�Y��)DhH�9����~
$G��5�ZP����5�,}��r����j(�e�A���-]���E�7�9� `hi��p�+4iY�4���\�w��6>9���@s�.���|{����o[���M�Y�E�N�sK'.�c�ȹ^}�7/c��/��7��G{ ]�|�z{����y1��Fmْ��s�6Wp?���SN����8RJ���;��x��"��^��zp	E��&�k����㫛6=n'��Q�  Iԝ?6e��
o��+��	�V� ��!������+^��g�@�cA��Dt��3ͭd��1��s��`},IA�����;���nd53g��&�R�c<� :�,���{#<����^S���XF� ��^��cnH���J�f�zbI���z����FV§�,ٵI�Z�ɾ2'Tp�����xF�M{?aɲ�~��oM�=̓�H��MP4��BL��t�������[�P\�Z����˿��EO)O��}��=��ԭ�uĞ���C���ڱǮ��kץgٲ�RSHG��/������?��O�|9�c�Gy��]s�=����L{K�]�¿Y��I��o��>�����b=�١���1�oƴq�&���O�p�|�^m^�
����GP\w�u�pp�	��A��c�wdg7�e���)��i�,Y�9FPJ����`+�+�N�U�Gʇ��U%�c^�6wL ����v�9��>�����=|c��{��v�c>�l���";e�J���,�Z���w��$�̂�N.�'y%����+��!��'��K���=�c�-s��R�J�����h�t\XK�����+�}��;�<��_�U���߁��xd�>�{�;����Xc�'Ň	�Ï�pX:��k}�<���#�<˕����ֻ��kiM4m��U��bMD�g�߳k�E/�{�RK��N�/��/fN�&βɫU��M��L<15Tw#�*���~�!*7��]�C?��ُ������U�)������o~�uW6�V|x	��M�yC�K(F�����G e�g�}U��0�!�!(F8�KxpN>ˉs����j� ��x&h15��"ry-}R|�+X�E]P��-���پ!�)}���\��,K�VYe`iV��<@\*W���=͖F��e{���k���L^t0��̋�5�I���l`pvڵM��Gg<%2�.��b�l��̅�#HX��G�I[X�R�j�����x.�:�H�7�CN�����d-M�-}O�^�ٞeH�B�]�¿ԍ��*����X�: ����g7�p'����崨�_ZN�C�)�Sw�Kբ��Ұ�y�L=�gV��63������{��`�j�� ��m���C�6�K6Y���ñ��?��O��uϐU-Z]�dp�^�7��ω�zXj��y�!�����*՟s�z,�qy��g	l��ܛ�N�.���k�\�"8�S2��jȒ�a�wZ}����R^A���t:o١���cɫ~����d�[�:hO<��Tyi�HR,��Z�]���\�YO$܋�U��F�9w{�x���퓶eێ,�ײd��h�;7Hs)��%�!N<�g�<���c����ەQ���	JY���+�{/�rqT�Ȓe��z��}�6[�r�mٱ����X��?MvO�<�Mأ�<��Q�O�Y}hZ��41#Vo���I�Q�vȊ[�{ܶl��欳�*�Rzy*�Y,,=6���h�(h�U��%�����C�YA�K/����R�S~A�?C�y��emɲV�%����0�����<G)��ȸ��T4N�:k
1���m�g!l����E0Od�Ha�}����׾6S@�v{S���ط��9$3U���-��cTbw����{�/�R��ozf��6����$,���t/O��q��$�К�q����K�+��4�7���j'�u*���i%H�^�mS3�k_��~����!��!�0(š����S	���^����d��x\�5�j������������gmbr�ο�,[vH2PmԞ���m����M�:)�4�?����W�>�,b��|�N8~��%����`��w�m~v�'bd1�J	����$�e�~�!�iXlR�{UeѼ���׼�5E/-"ea�qם�����w�/���b���nk�^�\�1cFA�Nn~dIȃY�A�J��>:���]*��f�!Ų!�.�Z�*8'�qxZS|E �q~��
���.���u��攋��4#�gF�TBV�ٰFS �j*F�ߔ���>�{d���`�Y�9��\��_~V�� u�/��H��V 1�+��d�`(�����v�/���7���������=H&�u�]^:f�-v���m�s������� O�֬]jûFl鲕����;�زQ{�)'y�J�����{�"ٞ�w�V�|`
���/�������ڹ��V�X�A��?�v�x��ȳ��5�竖���O{�����t����n!)���f�����G�f�����ۋE<:8vHX��M�9<2���Z�I��Z����I�߼�< ,��2�ʊ%H1��t}X���Y7���i���~,�s�<M���m
�CP�9�
�P6 K���R!���� �(2V�q��hgҔ؞`��d�QnA0L��GP6��J���������B��[@!R:3ɽr� �m\ż�H���Y��{��
 ���y��fB��Տ��Gp�q��e�t�HoH�߿�6=�ɦ&F��Y5�Om�dK�bkWeW\v^:~m�%{��-�u�D��c��V���0�)�΃�~�;��;���68�o�#%;��b��m�=�̟&�1�S;����/��ի�M07�ζ�~���{��%�\�A ��x�^np�7���H��3�����CPV0�1�X*���rW�f;�uZ���`I#�# �sqNA>���'��Pք���
^T^�M�`
�F�c|�-�׃����HB�\^zd�]�Cu��$�"b4��HT5U��,����e��T:�j�2ku�Y�	b��
���\��_��@��h͕ 17����+#����}
멼6�!�Q̳�#5d�w��;~�*k��ǜh��%v����Ș=��öb�!�b�Jמ�^t�u�zOv���w�{]R��ҵ``�|X��?���ߦ�\���j؏�3_�o|��m�в���^}�v�k^�Y�XC�w+gk�0, ������X�:��l@(�#��f0-66�~i�}pt�hl`6�\|��W�R�� ���H��Њx�b%|q.� C���C�V�`����Q�]���cbd��^QQ1B���׃�y{H1Q�2��}��z�R�S
��5������x��&-�
�ߖ��
�>]h7m�׳�Sn��f��?�{�
Q��r� �4�����9�������x�}~��󁒅�)
hdW)��*����y���=j+Vn������7$I']���G���F���/����v�=^�F��}�.~��*���MF�ʕ�=SʉA�����ܶ���.��O~I�*��<0�ԅ���pM�5��޻��	"�N�j2�l(�?�я��� Y���{.��U�����V7�F��o}�L��_�Ln�R0@��ɳֹ�{�O��;b���� ,tq��W�0G(`�5BT� %֮����`ۇ�r�b&�cP\��(^��W�ҹ�%%a�V?�60���<R�5@���D����Kmf0�C@y=�v\K���;�tx)�������f}�|�H�-r �=���Tn�09<(]�9�F~^$L);/�9^��o;���]l�Y�k�C������u#6�d��عծ��Z��G7gl�ь-V��3�X�¿�h:elddgf���&�s��o?��v{��G�\
�أ�v�N�e$�fvo��6{���{,�F�SD�����?�C��h������KH0x������_��p�YXjxp,�P�U��SO=5#t����'�E#�폘?CBRyZ��Ǆ)�}h�cP] �t>����G���,�I�F�JHIgA������>Q,JTV��;:��l�{�<���e ;���ؙ?�Y��Z���]�ᡒ��l��{��b|y�f?.|N�X�>�6bM$����I�p>���"���gV�����x��<w��7��	���o�=���u��?~��vc�ݲ�5��!�n����o۾��ȕ(��G���4�����7�X�¿U�N�ECg���W+W������2͎����h��@ڠ�b�U�z@ic0�X]*��q��;������)AE`"(������2 8�`a������M&�Q���+P+H�y��3��$P	�ך`�F0 x���q|��W0v�S+�22��Jb�7V������J̍TO�Ž3��4�P�PD=�{�k��_�F���t�l<��P*,��&� �C� g��A��R#h9{�����,���m�pD~�1��1xy��{���+	�������A����	ni�3��k_��?+�Eo՘nb��ݶcǮ�HH߅g�{x��T�̳Ƣ��GZ�Su���H��#ɵ���0=�:����i4������d�Q.��=���ܥF��D��44�����C��O��Ii0�0��#���M��N�'V��KL@��|�`�`�tB[X�k�軕���=�ǜ	A&*��?����x\k�vQ/���:��(�I�3ޟ(��B&+�*�C,��;dH �r�:����J9w
�%�Z>
�b����l���P�]�>?��`l���<���i6
%��(XS�\�6��9y/���l�|9+�9W2W��Ox6q9�}��H�s�4ʘ+Z"��K1���z`�(N
7�����=�����q��栘�A���G����"T��0XC��Qʆ�c+}e9S=�S��J��l�����d�Q|�+��E���z��ڸ����"b��lŅ"�7�\��K�D���E����BK�Pcq2Q�|sV�s:�>�wxE
^
�%h�������l��#��m(kz	d+�h���E�b09���e�k>�<�%)��ȥ㣱 ����ܷ�T�,�u�NA���	���me4�y_��tEPˍ�z1z���3V#.�>/�@7�̸�*<s*�:-�ޚv]{;b�yUڧĀ����@�����1��`��=�{�̣R����{��E/�{|go=���:Ӛ��6��?�y���aU��� �������>p�c[m4-�H-�9��mp�Z��d��ǾЖ�(��k�z�k#d�=�Ȣ�A���	�U�G-9x�U�E�by���Cשu��v�ɳ�x�X-�	%Pe���B��!ڦbU�������*��"�\D�z2��s9�`�}�&���aȋ�E�m�Iq�kjgHO�=���sYM����ڰg)�c�՜^uS�o��ٵ�bn�*Y���y���g3��s���]3g�*F�gV���_��{4g��sE�\Q��C@������r6�,G~�{�.J^l�.�@�p�v��mp>��N(`(��B`b�r���c"�Y�);ݫ��7�����b��u������0�O|�^�G���m.���:�_��`4����r�3zF������3|�*��8A8�Y�4AN�֕
�EA$�&!��w�N~9,�}ҋ�O<+hܫ��")
	J�U�b�n�2%1��IyZ���htXx����{�}�D͌*]��_aD�b��wQ?�)�U`����^������(�p�	�qi�,��YQ��ͭ@��T6%���*�Å`.�bC��Ҩ'X����õ��׮T�,��χ�/Z�P���8��hY*Q}%��g(�B0	�/���S���΋*M�0�CL��9kPP�2�uY������Py�����0�C�`�x�:��T`�)I{gEC��P�Vre�r$�cs)<�K���>JvblԿ��#��ƾ�[�x��5��PW�\�}�'�۾랻3je���3��"�.���yD�;����l��!o�y���G/�f�8��6�bD���m�շSC�J�Q�`�K	6Zp��TS�H6�m����h������X��}uǠ����Z����9����{#���|
�	�ݟ�{�C�A@$zqR"�^),	�s�~�o5fU�k@h��#HBВbGz�N��ۇ���w_	y1�$�4���nCumtm�l��~V�.�1R#���l�[]���%̹�Q���L+y�*q+�F2���^�c����X�¿���L?�g�5�.�Y��̔�� WPM�{��e9�/�_~Yb����f=��n�%��X�,/p�a�~-��u���L��r�|׎�UU�.s��9O�%Bϟ �,8��g�u�c�	�^��ye5*CT8�����$o	+��V6��:�X&b�ț��8ߍU�^��"�7]�O�S�A��P�N���X�VJ���,"�:���n�R�i/��k428�k5g�Y�	���3�� �C����V��a|1�C���ǿ�س��L	�1��o�/{�m[3=���L��5���Fĕf�`�j�ֺ,5Yڰlq�%P}��zo�XbX�.��r�^
v�M�0�F�L���k�cD�������� Ās'�R����}|��T�-*{�C�,oi#{GX3��n��_�ñ�,)�5)%� Vf0�ٯ��
Q��x��̫n�W�)�:8/�'�*,~h��>�=�r�6���a���O#�Ә��i�hOkϪ+\�w]�n�gX��sؓs�\ا��nf��T(ɐM�H�|�g`��|�X��h�S��j�K�F�/��P.qt�5�����V[xE����,#]�R� ��\ӔM��H@ĎO�4v��=]C'��=Yt�0�|C|�j�p����eD;��g��֊���1�1� n�Ź8V5���9��5[��,~,v?�FLYE ��T�?*w5v���X�3i���"���nR�P �:c�X������in����U��e�4��_�1�O�gQ.�Oĩ��L��֥�2
}]���u龳}���~n�Cy>�d���6�!��"_ �����@E�^���}(�P�fV�X����f�)�x�q'dV�Ĥ�G�mٚg�V����%�!+�����Z�F
c''��-vX�q�j�+`k�hQw~N���3a�^�NX�ҧ�PbP�G���GB!2g����PB�y��+K�90����a%_͵ܶ�έ��3W醨�Y#@�
��<�	U�Gx2��O��ד>��se�F>�=q�W\qEf�4��`�S������z) )�+�9w�~�扌d 73A��׭�ViZޅ�����K���~R�=8_�z���'��1���^�-҃Y'�p�y��g��@V�i��K�����
`��V�'C�4��7N5	��1�:'/y�K���3���)�:�&��d�y���'K^�	.&.��O>�j��~{��fcSD
!�[����`Y1�Ŭͤ���)dU����GL#Y��F���QK�G&	#*3)C	����!O#&��߅V 
�I�<"�F�Ne�
��^P"�G�\
E]��1>7�^BZ��V�̺&���:G������JT��!��2�״6���:�����9���z
ȫ%�Kq�n�[�Qݓ�Kk�כ-���u�s��j�+�"3$�5�2���G��^��N8�=ϥK�����n_?��Ńv������lyY�9�t>p3|���U�gVOQOG����|�7\��H�HL��f��V��&k��u�i��op��L:�~��~�7��_���\i\{���]Dlu&�Lc�4{�N7d�kX��%������Ɋ��YC����Z�Ŏ����N��ڬ�.��(����u-<�d������,AS���z��u%���6��/(2zCR���o��0^BK]���u�μ�V�iD���T�UDl����Dh'Z�b��we�f���lC��O����~ �uZ��W��(���!&���d`R���3�p�oȕv53��9�l����䦧�_�G7 �U"�P	t_Ǣ�y	�YI!�Ed�j|/��"��񤝫e\�qۼ#�j�e98X�ɴAN9�$[�f�O�����ª�P��K�����|�7ۿ��������^�Sة�	Pa�sI�P	C_MA�� ���1K! ^��C�G�j)���'�
�ٯ�r�3v��,x���_��(���Θ��/
�s�]�ys�L��zI ꘨e`Ȼ�=d#D�s�L*Qu�����y]�	����n/?�ZPRН���Q�1`�ƺ֩F����Y�KAc=��&
\x5Z����4��a��⾋Ɣ<���Ø@���կ����J¨lN��(�8͂$���ڵӖ,�����>�[�/|�Kɀ�ϖ-Yj��#��q_Ǣ������˽�����^��+��9�H���n���Y�W�\�=8O?�,��<X)Z+^�	D)<��#>���_����|�#^��f,���� ?�5��׆CyQ%/C�v(�'�9��~�(9~t/j΢���5����lV,,e��������Q�Œ��$ "�����qi.��z�h�Ȑ0��=�/Z�<�JR�1�'��R*�������R��bs�H�t��Z�E%�EZ�s��'[U+E�YJ^�+���q�6"�罠���@m�7%�̟����c�~�^ӱm<\0��z��ב��нy	���0������R���7�>	~��~��6nz�n�����;}n���=�<[��P'�,Y:h�~���_����^��A��v[�¿Ճ�59Q�`��]#v�1G����d}�U�?�arٶ�q��Yv
��/�ݞ|�q;�e�Y��RW_|�G5jg!bI���p!I����ۇ?�a{����3ZGmj�|�6��(l�}"@X�����k\�h�	o]�g��9Z�q=>��X�jT@�8�\	&Q��[B^TG0N~7z�Xx��6*�X/E����xu�*1���u�־p`�S�]T�A�-���y=Blj���C�3&�˜0W�a���=�X�ū 2ǣ�E!U��FC�q�Z�_/��@�+��(
���e�����'wq-Y���;�1��3'W"(��<m۶=�s�C�����h��=�y�k�A%��g��w���2I {n�3v˭?���m鐕�%{��_�5�����^w���V��UW������vNI��Ƣ����dc��\ȍ��N��m|�Qk�ǒ��O�t�UrL��o�޴�׶l��w��}�ݑ D�M(�#��F�W4<�dY�
|F7�׈L�N�!��M��T�b�Y���М�sa��@8F��x��
�,S�	�X$���*!#Ꟛ���D�I�="^�Z�RFX��	<:���l7�' K[ޒ���.��_�3w�F���������q��3��U0a���jq]��՝{���7�!�-4�5�>��Ϻ��� �8���q��<��Ig������ܙ�+�?�
�zQE�������o�o�q���\��1��?�>�[�y=��Rԭ�1{v�S�s�6[���zkmbr��Z��}�����ˮx��AA�u�v��?rJ�/�K�3&��Y�kIz��^nL$��u߽ގ>v��o8̞����L�?ɽ��)�oO�J��Э?�Ņ��ظ��8{j㦢 ����)�.���B�_����n�tz	8Q��^GFE�5�G�g)XJ��\��,>5���*����BB%$T�����e&�@4Eᘂn�#��`�ApR�k��vX��/4癝3ǡ����i�iw&�u+w���Y�\�փ:o���v*�^�J=(ʔ�����&R�������|�yWp;��el(�4>9QԧaD�c�F��@�ր��+Z���״�bn���]�J��v:xql�O!�F�<CFRr����oذ�~�#u���o*�;��Uo}�-Zb_��W=��o
k�b�z�+���+�mz�qk��؉돰'7>��~��F&_���-�����V;�S�_���Jo��hvx��@�������;��;�V�\�&��I_���u�G���6�`�)X�� [��1�,(K���kXO?���@*��𖷼�q>�,����?m?���E@/�ᴐz�N�Yt�8{W���B� ��,�����o˞��>�@R���^�Ғ��+!
S�uH�I���|�>�];-���k�gAO,�p�^Z�zL�L�Z�+��|�[���gd�Ǻ2���	B�������&6̹+�r�5��	2�ٹƤf*lV.5�&�������A��KVt	k_�����s�X�b)
����?���Z+���~��N㦮����<�����{ϝ��C�@J@�S@E�����T� ƭ�2h��� qd�	':DM< ��g6�A��+Ib��v�����R�d�?��S��-�m�&3�Y�T�R���L��h7�@X
Fbc��	�b�}�;�q� |�w�w��?�)��Ul ыJ7pd��������H�0J���	�$�)��<�J����ıD#J���P��I��@4��D.��1"�U�
���+���������;Q���>fbGVH�̙�ye�:� �ǅ�G9K�k��(
�v>g����g�W+X'*9-�W���fce־_���ݳ�{+�L�]O��:��ÿć~x��n��!��e�ā~YGxyt��|k�����m���y�!i�ҟ���N��O�s��=���o��VK�x]�\Ǣ��L_���0D��rˊ��Ov�����I�*-��!��X�C8��t�y�{�:��ƥ�'-ߨ�N]{�L��@Y�)��ׁ���
03x��4���V=�$P�(�)I	+}w��kr���B�\��b�;RW�rHiʒ�	Uz��+��>���6��ˡ5֔<��{���k� �
d���?� /�Y�����%����,�)gP� a�
���Q.�z9Nީ�J�=�L[6� �`���c��BI,��3�bє�u�O>n�F,@�%�� �D���-PE��O�S��4��i}Y����<:�ÿ������OL+s�)�ۈ����i�>����l��z�ȏ9f��t#�+K"�L���db}9������H�Q�H���l �"�;�3N����Z�!��|���ǚ�lv�HmhY�F��1�����Y��7R�$@�����R�n�SѱN��G^�8�ԘG!J�1����������6S�������P�q�ְU���yMA^�Q�C8��"��d2�R�z�/(���oֺ�ː�I�����?��X�)L)��-TF�c���$���O�q���-�׫^~�S�K��p��ۿ�A�w���M��w�y������>�o�!���[Cs��_s!�m՛S6���Z��rr �ג���2���Ĩ�5�!f��9�E/�ͺ�wgg3`~�a�j�a�;�OѶZ�VV����Ln��'m�ݾ!�p�$&M�*�t~YbJ�<� �"ZR���lC�����`���q 1��6	l,D-N����q�����=���c�^��V]A��y��"�^����%mJ1pH���+Ȅ��f������^�g.�_�M=7��
ݕ��uQ2���Aq��0ψ��=A2~e�j]�X��o8Ya{�F#�k����xĠ�����i�=͵�Ѿ�Rkv�L���mHc��{�s���W�ʧ���8X~�m���<;�XO��������X�3C�������,����lt��ɦ�|��>gcim�Tdh�
�&E2�\�¿٣����l���^y�����s^�lOۮ��l�����F�(��Z�R[����a[w�R��#I�[�8�2�#�KO,�E1(
�ن,���`U�W�_�;���}T���X���r��bPL�t�$KV�
���A��C�Kx�*����v�������n�M*�D�LP������υ�h��f=��1��
��2�A�1j )���`p>QL���QS�L�Ab�b���s����]��cnj��r�v�ry�z��0�-�=�N�n1�00�{���!}�!;�%��3���۞�F�φ��:��4�v�I�أ�lLϻ�pF_2F�3��w�O�&����;��9�i��g.8��$�WZ�@5�W#���:�t�?�g�Ɇsp)�v��.*0m&���l0�?��?م^XP�b���G{���ͯ`�\��%p�0�YE���>��f�9����H��s(���C�0F֢��V\��͓!�\�AyX/�>�5<��"��h���6?���$%X��P�e�� �,ƙ���A����H!w
"�Oтǻ�F��Z;����C���ľ�,��̚��o��33��o�s��&�^�9��3��潔@l���-oՍ��z�a)~�'��7���>��[�;e0�&Ӽ�\u��ܽ+}~�m����J�犲�f�d�Ye�^v�{�z�<{�F�����/�Z����'�BIf�;��~�n��&��5�Nx��:f�/͝���'7�3<n�rՎ8�(;��uv�y'���MǺb�p��^z�M7��"�gS1�K��B8W���Eb)0���lB9&����|�7C��K��{D����uQ�-o"R�Ua�XH1��x��l�wO O-��cEHE�L	��6��Y�M���3R��m	r��P�;��g�a�8����D&�����W1�"~��dp>�����`�2�*�9���i���b^�_s=)�Z����z^ܭ4͢oN���\���zT��*ʹ���
쿈�NRӿ�����\�h�����/
�ꫯ����ﴖ�<;��+��,	�I[��4۹}�y�i72��ɲ">s\20/����~�	�������n�G~�ȍ�t�N���*�¿�G�Y0Z��ot,���K�y�?�X{��׻u����/�ڵ�rNu�l�L�S����X�r�� ���o���_��c�4��;X߸���o��"�3\�cb�	A+,D0bY��,�IٿwW����/���<#a؂��6�%Z$�*�~�И����?
��Y�<�'��7T3ch�ƫ��x��3mB�<X���_u��.R�,e�
�g�x�j��8֥�-1+���3��^�?�x�.�����Ox�bŚFsabE���B��B�%��J���L�dk[sR}�ݾG�K��BŖF+�q�Y){���m���Sݽ�^^����~eE�&`�}�_�ߏS�eyƬk%H*7C�c�Ĺ�/�ܾ��>�ev�y/�����)o��x����������lȊ�ױ�/�>�wı��Ѧ��g>�Y����� �v�����8*���6:Fᬺm߾���o�օ��ZL�����x���������.� ѧ>�)_���]��ψPL��Ŧ������ fHH��8� A�(PX��s��糲U�AHΏb�R���
���:�%���M���D�,T�AX�|��2�D%�
�1)�z��_��_�k/%ſ*PƘ�k-v��Ǫu�kS��
�	$�.a�3D)�9X�Ϫ�C�T�����JaP���_��`!�i��>A�F�!���"��`��H��9�%T�NtL�@5��`�:�t�&.������d��Y�ֱ��ã��̳ٺ�r���2�;STޑ�zŹx�=O����\��x�rX �7q�o��^%��K.��Q�s�)g�`�LN��̵>�����{F��j�k��V��_Gg@�QY����W�CP_p�Ey�⩂~���?�1woQ�E4K9Y0X����Q�෾�-�.��B/�@�@��
D�E��3,y0,BY�
؉��*E	E�D�Q�/����|��F��.=��r�=�C�"����@
�r��'b�,4��7j̑� L@����ΪT�EtI��Z�ipN�s�)���2�J��9�[��*!+[qU�d�c+P��c��cL`�!E�ʶܻ����c���x/�"&҈�(�]p~��'ltx�=���6�kGz�n�[��R�"@#W�<�,�Q돷#�8�cqO'��^zzs�-͗,�93�=�,�'��X����Po��@�-�l1��s�v�w��x��_�m���a�g񙆓���k�X��sN��?�Yͥ��q��/u���d��M�\饎�e�Ъm|j�mݶݾ���x���k4�%0>�Sݙ�����
�J(�E#�x��21�*( b��JP0*-�6�'˓E�LD%)H(]TQ����'�������#��Y"A�� )$��n���V(�eM�_�X�!���w�k�Ϝ��{|���3a�#`e�G�q���C�Q"�N����wz%��x��ށ��4Шp����5�Dzyg�\u}�A�ɱQ+7�WI�F_��+�Y�MU�-�D���X�]J
#c�4�mE��h�s)�/+�s~��l��r�AG�^�L���y��
2�JwH���o�F�G���xR����p���y*s��N�j#���x����e��RT�^�+YU$`d�{˃+�mg�wʭd�!�x��;�g�UC�e�C�^u�U�(O;�4�H���T���&�5r���| )��X�vK�ɢs#���d��'���|*=��Q�?�ѹ7�AX��? �]V��V�zY��k�J�Z�~��`���)� L^������)oa��TyS��UDN�[q<[�?XW*/�h�9��b�sC(���'��@&�kdl���wHA�
*l���E���~4�C�.���%i�٤��[�}W�fΓ���̠R��M���ʜ���{ �v����6��=���J@g>�|�W�*&�{docpѷ� �bzzf�ڱ?y��2�3Y�6=�%�S�!����݋�S{h�sT���g.̸R�t`Z��m�ˈuWD�t�%�_�k�� ���`���`�F<�k`�I������E���'?�Iߔ�A�p��?~-W,�����W�v&�)���,PY���c��|4�N� ת�c���`�^\R�����p�E�YpLE�8�0Q#m�K s�Yo�f��|.�iމw���L#�de%�u��iK��ol�+v�0�N\~=o�yQ�D�7oRק����T�X��x����p�u�0o��$�T�GU,X�s�%�e��X7F��l ��{s[�)7�j�	�d�I�yyh��@溪bB�AmdD�����y}��_�}N�7���������̟�nȐf��J_�&��V�Oϴ�ɣ��~�ûlp(y����ʔ 6��F�$���&K���6Z�"�~�E���f��d��m�z���K�1���R&,����� e! (���O���-n�IH�d��h�h}Ja��#��%oɲT0W�Q�'z�+�:f�"�x�AB���E� �K����0R�N�
��F0�@�R�Q)1
Aל�ZKi)�b&���<������H�a0�7��%�5=	 ֔�y�����l#�1⻕�a�r���I!���g#�-r���X\�ۂ�Ӝ�f�Y�i�%%�%~a�;%t2p}U��t~�Ԫ��!*�8�W^��ɑ<!ŋX׼Ϗg�潒�HX@`��dՍ��'m`{��J�V�Z���I(Zg2L���Қ�� ��}5�x���du��Cm�ܵ,{i��H��Rő4��0�O����[9_p�^��w�>������M�{d�S�c�,�����˳keMŠ��T HG�B��x��rs�Yd[%�D�dh�r܇(�x*׀`'\�d�q�QF��D��7�hΫz4�.bYDG*cy��[FgPS��C}�f�u3�ۿ��΍����s����<+�*q� ����ׯ/�S�]�j��bs
&� �G��<)��R"XΚq6K~OJ��[�E\ks�,b,"Χ��2�ߨ߇ ���N�C�VL��<MQm�3�۩�1���<��|��6F��~��Y�H}���+�$x�PQ��<��QfK���0�־A��\��G^�d��3{�g���y������_,�i*��^|��2�a����^_0L',"�}ڵ�r������z,��c�,LYw�?`���>���x�*� �BP����[��#�&��,J���Hu�`�}�m�y�G�x�l��1"J�P̭�%�n���@���8V����͛zK��,TxO��I�L��Qָ�4t����Cl.�A�~���$�8�g*�=�f#)����ߏP�{E�¸)&#o&��ϕ���܇��R�ϲ���D�p~]��}���o~ӫ���?�q��C?���eĐ��׬C�劯!�F�}��1z����ح�0�j@��EL9��큪�k���/��/�ܲC��h���;d9��Դ���zt�&�F<9v������mL�(j�oh��Q�H���΋�#.f�
��&P�Y׫�$�#g_�X�F�'���{���s&�G���*X-���P�^��+Y[H��!K�&^��Y�xK(�X�ZZ��-?x(O�q*)A^S�G,I0SPV����-Ԑ��<f�S4�͖�"���ͽ���*�`����-'k�Y�y��5���%zp{��kDa��%(��vT�Z�>�`1����6<�*��Zӕ���j�i,k��f2�H���HY��}/�r`F��e){������Y<\�@PDw�!�u^4%ܦg��R�����9GW<ZȲ��Q��b���$���~���K(�]�ML:k��_���;��$�:�[c�}_�sӼ�p��7�SA���@y�E���yw>/A"��WF�^cJTQi���s�j:�֞����4�߹���ӳ�wLcy%�G�n=�z#=���*"��6K�P�-*W�,�w�`�����<:��)���Bs~���x��PL��D�P��zS��s�[ƙ���dzɍ�"�n�1�:iN��|��¿���5���6y�	(հ�ZY<�'�]�/��z����fV�g�D	�J�m1���[�i"�:V,�SP�S��'���}ˊτW5�κ?1o�㗒yH�JTN��,��Y�m����ڟ�=�OV���b���)�d1���O|��1�S<��D�%�y���He��;��G'$ة����^�������b�u�T��'w`b�&Y��$k�{�f]�X_{&y1��z#�1�ǲ� � ��ڂ�<�k��;h>y�R��baC`��@�xn������9�Cc/0�����F/2����,��=���X�¿�m�6��$,�k?:U��m¶թ��6Fw�7c\0b�t
�ο�ń�4�C����F^�������5�f�ĲuQ�IE���_�F+��F�ә{=�,�Ҷ�ע��:b#��<���&�'���a�#�FU�-�!VL�W��(/NTP�(����� ����wu
���9у/L� d��Ne;�!ť� \1��S6����,߱d=[s2��	�	/�W�Z�!�\[�j�-]�̃��t<����.�O��ؒ�����Plѧ�*%�h�id�Ǖ8D��g0t��)���d�������`�9`���E�pl������/{���DV�m鲥>�Ln?cc�6�d���Es���
�B6�Ц-0�N�W>.Ta�L	�t���(�'�vۣIVP�s�⎐N���Y�A�N��Xݓ����+u!GTz��Fe�n��4���M"B�����.��~XX�w8�o�D��9����w���{^ÇzD�b�������\���y]kGA�R��	r�	�ס:R
x�� 
 S���p����jVճ����o��=�P�m�>b�G��i�
��*�G������|Kqʛ�BVv;����$����iLi������u�o$'��%�<1��o��\����y��'-+����ױ�k�n���vZ��	(}�}�km��徙֮]�Ʀ���f��[�~��<-	�G6&�@�տqkK�D���f�p����v�
���`m���i���xq(����"�9"]0ޓ���y�qn�:���v��y�}����O�J�"�M�﨣��F��w�^��~�Cr��,?������sX��\s��7��M��W����_��_�b@���}��zPԮ!�Tɂ�����*�G������5RD��5�C�9+�	��O@�G]޴v��p��,�JF��9y�q���=mKl�r[Z���J��)����$���MO�j=�G=��b?�'Avj�Ɉ,��
�F�q�Y���>���m��?X��%Mf�_�'�hc��?Psh��j7��ױ�?��f7�VGI���s��n^��Wم���d�(�sءk�g��)�'�z�]w�u�%�41��o����o61�෽�mnݱX���/yIg5[S@uY�>_��~�~7!*7�xV��18�4|-v�K���������{ /�	9�����VR�o,�D�����:2	d����C� k-��ɉiMTp�D�Ku�ԴE��=^\$ŦGy�8< 	Ш���5����E����iT��?���(�����n�����.U2�%�Ջ��:5s��U���k�:L�\y�u���-�\��ǾZ��w�@~����,bE|�w��C=���_b�]�^�EJ�ܛo�E��=���v]�����l��n[~��=�ȝ�>�~ g�v��=`䙝Y��$�)u�[�f�x�Ŷ|�R�ԎO��&=�ӯ[Ln��I8�����#�����޸%R����]�S���?���`_��ל��~�Wx!1<	Tc1<R+ƓO>�/�>�����3���ҏ
����	��Q����+�O�����;����R��I ���תe���Tc6���j,��CQ����Vj/����}vֲ���l���:)q<��K(&��}}.*o)J�n���uia=�n��s��݉-��-�J:n~l�^_�)k�WD��9�6�VS���8i����������#��j����'�3��ח��d8��H���E��e�'�,Kط<�E/�K=`�r��V�q71:n�sn�'}�L=�ܳ������m��<kU:yy��zꙶ����C׮�+��F�=��;��IF���>�9��N��3N;���^{��Ǽ\0�T�+����\d*�L��)���,J��~�}��fk6�Q)���
�"I��Ijg�3Z��<�x�#6.n~6�m4Y�p�I�X,�o|cZ���
.��`��Nq�9)g%�}�"svr<���z�Q�����VI����}���I�ޣ3���l\��{t,�4~?�WJ�)�K�)��g�3������͘k�ǈ��ێ��Ȭs�w��y�������q��z������V��hbZ�d�o�fO<�m۲�1�ի��I'��%����)��d���a���g��c�G@{��V���\�d�Vl��ەW��IcjĞM����~b?�$ؓ�54�'|��m����9�BW e,e5ؖŀ�Ǌ�aA�z�E ��&j��I��5im�[^�="_XV�g�Q��6�P;:�Pu2p4�	ୈ�a��4��HG���y�+/A�wI��r(Ы2\ץ��=<)���p_L��1�O�ڪ���;h�e��[bj����b��mt���^�!Gk�!��������M�~��ݓ���^
ts�>^�k^�;��#lb|��Fw�/��~�������l	r&I����y�A;����QGW���w������.��|��>ϑκ�c�+u����Sq���g����u62�ê��my��$䟱�]f}G��� ��:"�w�����9�W��J������g�E��br�>��F����{�x���}���*���;�Y����k�+�$'a��6T�+6c���덂Q���*9��-��_��L�+����P�G���"��9aD�"���1^2�2���|�
�1��n���(���X]���2�w�����GM}�za�0x�r���w��&���3s���gG)q�?�"Y�q._����*▍���g�d)_�k�8��f N�y�+_�kO_y����?�coV�o�Ϳ�?��?񹈙����?:6l����Ϟ��H��#���Y�i�9�A�뮿�N=�,;�����Î�N8�6w��	!���;ow�!����j'�t����X5�?��F[�jȎ?�����4�c��J�W�1۾c��%�Ɗ�k�a"�ُ% ������C�1���C#0\�ˢo�34]��t�c�AZm']��Ϊ����<*���������Z�^fA�H����6��"]K�������X�y	��>/ap����e0ڨ�
}�=�s�;���E��k@��;�����;�)ԧ e��4's����#C�f�3	o�S�����\�����^c��#���:�,�����!u�t�MN � 6��u~�9�V�f?l�=ro�)[�n��?��F�G}O��Q����ϭ6<2a?���X�'�֭q"
��=�Yi�y�^��X��d��v�y��iR[^5���n�7��r[��{k���"ob�N�ɢ�8E�Jε���<xKa-�9����*ңW�EQ,7���p8a�ެ��Xp���ٽ�����}s�M0:��3����R@ΌH���Y݆�U��N�������)�/�P���ΊMlP�*��y��*�8��ň���ǡ��ӈ5�E��#�TВ�'�C��b{	�={�uf
 �N9[ڿ�S$�u�?�;�:����)��X�|'xM`�[�pσܗd�2[�z�M���FQ�u/�����a�Q�u�s���`��w�{lx���v���E�����w!\��g�ޘ��ݝ}�����NZ���`j4�=Ѣ\��-O=h#o��/��{׻��X�� Y X}�����z�j�k�GKMp��ǋ�'��%�c�_���V6�h�6#ŲS�+�+�!�XL���*�|����U�}a����0��RL���k�+Ll�Q�C
4�q%�s!.
���	�+r�9��I	h�u����B�뭲[�e{aÜ�q��}W_}�{��f���|�����ݣړ!�9�{��s�l������MM&�0>�{a��¬zg9���z��f��
�x¿xT{�����{��ղK�V��*�_�����¤���P�ȳ--���
�����eu���{�m_�e��K� "mADE�b�h���-&Q�����"��b�-�`��BD�FT�" ҋtv�������|��~�9��{������ܳ\�ַ>�yN���]�AY�x��%/	��������,���k��qՒQ�>N-��U.���f��Y�x-C�(N��9>�#_%��lk���bm�m��R�f}e=�l��g]D�)t��8�����|�]���g��X���/�:�|�Qh))JUH���<ήJz�ĸ�X��u v�׫�<某��c`YW��؅�[#��i�9~:xp�VdG�.}� �>�>ѧh>*l�e�;4`sk��q8�}����Ͻ�֮���2d���� ���zu)^���oV�':0X�n�`X�|��$�H1�É- �r����� �F-6��A�bn�\~�_X��$6�`}��Q֐�?Gǘ�^i�öYub[�2�═��Aơ8h 9.�Hʿ��|�X� (�FP�V��H|��{�j"��~А~���x���V����7|ܾ�8tͲB.tL�`g<LQ5�L��;5�,���h#[�<�s��ʿ���a��Yk�=eH���\�(��?�nr�c�Q�hw��.ŕyvg�5�7l�Du�n$���Y�/�"�����X��<�Jޑ�nl���۲�J�2�eO��)���wo���w�)ny6]�W�8�)���1�0��+R�ʩ�|�{ʽ)�#���I��O���]�7{�����E�Ѣ^5R7�L2X��e�s��$�|�IV���Qԋ�o�L{�4��e�����ްt�n�)8���kV?֬Ò�W�9�^����%�Cm�3<��6������������@ ^�e�h�Ǡ���/FȂV�2mi�T�b�J���bT�H@_!�H�Gh��RӾ&J|XM�Q�y�b�",�u���.�-PW�����`R����V=�Hx�I���Q9/���JX�t����[n�3t��y�Q�T��r�%��:�[�떱��X�^�[���7|���8&�tW�.�v�����~�oX*ЬZ��/n����Ï�vTN����7��Ƴ8w�q9}��3Xy�ќ�MqKK�e	ζ�egY��|$P���լ<��I��S��OsǗ�����>'*��������|�0��.�̌=��>��]tQd�6�o��݌qu���¦�=Hݑ��m Ϙ����;<�ȣ����]����"�2�z�O�4 |7��J�և��7G��~�3�mrg��w���M�{�N��`�5{n8ꨧ���=.,^�gN?@?OY���s����Y��E�j����7�y��=�4)ShK[���p����(#�Q�=��l�Դ--,�5����WD�8�a����m�<(�����%��P;$��u�3CT/a�=��fox������j�8��#�	+��:�ظ�u����?����R��"��dfZ��&an
��/*�+���85�}��ap�?�ߡa���	kW�
�7�7��yX򥳣'�^Eϓ*K�����0��2@��Q�*���}p{P�L�|M��a��2��4�k�TO��C�7����a�\���e3�o�6jz��Z���`�	ƭ�>V?�"���+W�Pm>�⇹_���I"�s�!����懧���s@��Ca�ڧ,��v�,�=�[�(���Y�B�7�䧡�ws�M�Im�����vا(��	�	��VC�˾���j�S��SN��˼��¬��aϐ��VK�x��|�;V��V���e��x��h�nv�@�ɏ~�c��a��Z�CP(�n��۲������M-��q}�-ʈ�K�N{�*�s�����{J��n��p�Yg����}�d��#�/E_@��
B'�+�/�z
�^t�������9+,�u�%�}�'�,�������_�첼��r$�-���E^�&���/̒QI5m���L����ζm蝑Z-�6eE_�r�e�a�k�+,_��W��>��O�M��T+�_��B��@��mT+����g>q�rN����ծ[���%�r���4�<��wɋhDR+	kO�,KO	6_il�`����%?��U�V@�?0ʒ�_.�x�ڟ���U��:0����y�v���(9��Q��Ch����E����?/��� ~��*DЧ0�{(���;�x���g��Hݠ}P��_�����|.�J�'�]ͳnf �:�R9>~�!�ED�o�`�P��}����eM��R��c}�N��4���~�㟲���^�|O��Ю���#��!%)k��MB��e,K��O�h\�"b��7�#̂��0�ꈕ�+6=d+
�}��TV�k�b-�����yN�f��G��U����
A���3���n+�&������O����?G_d�Ϫ�):��/���i2E�U��v�IR����i���f� �{O-"cf"�r�?�A]�=B�_��W�k����eFY�E�<?��,3\{�V�s��#?��T����f,�_�Ѷ����0��=���n��PTG���R��&��o��P7�6����yG��޻�W��+��s��i�Q��C�AT�°H	8 7S��$�E� ��J���ۙ%�dmx�6��-B@=�M~OG��X4"
�RĈ&����j�,OO�e�����h'���.ޞ"[���5LjI�GA����������&MGƃ����i���2N��E�k3kV�Q�Jɐ+i�r�r����W��($�y��mA96%w5�՜E0l��/�B�&�\��%�7���1�ph��~sK�H�:���>k�H>Č��j3�ᶞ��?U��9�����P����z:�j)q[�,�tp*$ �k�z�ue�{��&Fb�t��(�d7���<�y ��+�q�WGY�ry}�F��� =7�?��s��t��X��u�v�U#j
�� F�LDj���m�r����H,
o(t�SnO���UDcK�Y�'B҈:z2E���;�1����KII���@eT�o�q$�~�9�OCh5Q�0�<�@��H��QJ�s�/H�[� ���/�c�h/U�(s����z���������>���)���
���>M8;\Q�&WR�,��lT϶�,�� �b���k!�|�;��c-fċ��ѷ����',E��1���[�Z�|!J���X�s.B�t=4h�Y�:&Ÿ5���h��=T�������Gu�X�;���Sr���)���=S�xD�!�U�Y�IcE`_M>٢1�á$;���б+��ΈC��ԒQ�D��'��W�u�Um��)<�n~1��8 y�˅�Ȱ5��f�%BX%#�K�~���=X�J
�n��M��Dj��V�K�����?KWm�MT6��ь��U]����\��)�	�w�+m͗)�Q4ΙE^�p˾� �$at�W�}*iE�h{���qkI=e"��m&
/�2%�\��EMqT�Y+�;�[�PQ�Mݴ��L�z(sQR+�9ޘ��-诮k�/�m1f+�w���dS6{oᘸ�,TB� >�篙Oו,�&o��y�	�Q(��s��)�Сs�O�_����2gNOn�#D4��Bm7k#y4XN�Q�/��C�1�a�V�6h��e_�J=�7��Zr1�0)%P+��>?���)�jV�7W7��7V�Z�u����4T���|����{�M��=��1��n6�=)"OC�WT�Ÿ���0��l-�E*/�,�re�v�0٬ �os��$����>,�d<��Aw����U�E/�!�@��C��X ���/}I�m��ro��]}��Vs���dJ=��Ʈ���/�xw�dd�"R� �'bl���$2BX��x��DSH/��-�7.�o{z�,�P�s�m�W�(�]�R��!:�d�y%M�p�J�J0d��\�aK�A�����~�s��y=���<�տ�Y����@۰c��3���Ot	B<Ǹ$�c��p��Q����b�����n��-��1�T4��șlM�k�B8�evi�x|�+��T��RMR�w���B�#d��q�$�uHť�b}�"�h���Ȫ'�@� cJ�ʾA���d��>~��*̼�9����5�8���d+���IG�*�5�&���Ƣ΅��k1�$�ܟGQ|��������x�5؂8,�Kc0����馪[ �a�m
LʉU�1G;;���\(��P�\�|LZ���u�!�ƿ���Q)���l
AC��\JW쁡T)��;�)r�W.���(&��A��H�=�C���{p4����h������g<>��̍�&��8Z� P��j��eU�I�s
x9��;��H���9)t)r>�&�硲*���#
=�O���X�"ߏ���T�E&[��ĸ�CD��*��h�Z��
z��-T�̪/%#�Gڽ� 3J5����ǩ=V	��~��&��[����\�W�Q�y������5)Z��������aJ�T����E8��Uμkiv���~���7�@�����J��9�ƴ;�o+2��x�::+Yf�ìl� pߌ�;k� 7Tqq���F��7B?�Z#񿑞�ږb�����|%<^��5�h �M*���B�c�R��������H��EM��\�{�"�7����;�;O���;�֌R:;���x�o��!����iҎ����g�C���Pv�Vݛ��g���c��E�wnM�y0�chA�}�g&�����3W�N���ם����`�ީea+Bf�yXI5A}}t��2�s<a�i�����z�IM�3���L)[��m�H�T�)e0�5��"@
E�SL�m�_�BXF%�)�k�c��L��SD~x��d'���O�z�a���m"��V�7c�X�_罴����}K��z'��|��exoK�TA��[�mlb�ް��'=J�x�޷���ֽ�tY�=5��\�3�֊�(?'u���|�ӣ������ȡ�S��Q��T�F������Z�q�CU�$��y�Y3iy�!����o��Ψ����)nx޼���a�:KΤ��(aҹ����M��h�7JVB,������ ��/Z�>f_T�� ��%哽�8�9mmry[$O��J9W�G��U�x��=�x��<9-�x
1�Z��S�L�xX�{=�Z��S��)q�v��&)�V�I����"Aj�a���[�$)%�v��a���c�h1U�I�� 2\��&��h�VO�q�Q����PV璵��r��y����s-,M(��`s�V����:`�A�����,�ߕ�����p�QG��sS8]�\J�}~}˯��<��Us"J@M�y��3��{��lq Aʊ��_n0Pߔ��58<���@�b_֢�W96S`�|����~���� te�q}szYt�WŅu��3���
!�d���������d���־��V�1�R��� �c?��f�7���crkI��b���?����j�	��� �[��ih�/������B�Y/*����ہh��K)�)��;��}�1F�ĢE�æMBGg�l�y����52+J�X�K��a��/^b<�rw�m�d�v�a�����y�T�9�~��������o;��W�J��q���w���ۢ�"��|ޚ�R����)Z��f��Dy���yL�"�u�$W�����.Y��&�S<~"��H�z�/U���@D?,�e����{P��M��D����8/�4�y`��+�YN�o-��A��-��Uua7�l���x}QS�1T�e���3�����~�Zu+�
�y���c�1Ѐ�)��y�q����~��[r��$U/'�iXq�I3��Be�%K��A� ���AR��eɀ%{W�^c݆@[tvw�=�\�X�$�_0�������������{��^'�/pMn��_�j���Q"�R���/���(���b���=yWq���B�ޢ-�#��믿>�
����B0���U���+o#���xg��Gl�	��ҡb\�;�L��E��Uա��>g�y�s��1�W���>�_g�>���=��¶���q��?�����=蛡t J�����'>�<Q�y�E(���;#r���[��H�QI�D�澰ے]ü�¢Ż�����ʹw���R��k��^������J�ț^��4gx�s�-�y�TNK�~�âӢ��O{z�k�ea���V���f��C�A��.}<�ce��DV���6@��XZE_T~>\����mg�Z����?�c�¾Ta-*
�;-@=	r�P���*>?��#I4&fb��6�B�\���?F=lUU�f[%��,a τ���%����w-(|?��s�T�2?-����u��`h�m?~_%�Ѝ�������*��g?ks�¿׾���P�P?|򓟴�#T�ƴy<���#?�@'��=em��֭��"�i���Jٶɼ��l�΄�ǳ�O{��L�ɝ�g\�l�p�����&�|�/¯o��ݐY�������=�����p��Ǆ�p��X �|�t�bWEA�k���lٲ|" �JV�౎���'��mU�H�6����,l!���F��b�ɡ��呕�a��}�"=��������~-�o��|��0ط9��prȰ��Hj!-yL!��rHߏvr�c���g�����և/~����LY11��ΒmC���ů;���SO��:8���^���/��b[���7m;�9A�������@�>��G�7�����'���=��~����"�(�:!�C����|{z�V�a3^�w���`�شV���n��e(*�êU����-���a��e��]�f]�ߟ�8�\�.�}�����'[G/�w`аYYY����c� c(yؖ�+R��OwԶ�jR�*#�oB��;�p��z*�4�)������p%+�V�U#�z)q��0̖����]��C��ې0�1E8������'yY\~�������ֳ#�0.ޠ8���z�E
LCu0��ۻ�=��*�a�����Ɯ���S�ׇ˿�p�	��7d�'�n���p�]wY$b[��i���&E^p�E݃��|�����/¼��a߽w���#a��}��b��֮[���p�?	���ߔ; �fbrr� u#�+ĀO�]A�����}�(i+�)-�e���"�C�������~7S�s�N�<GOs`CV��5� �~��hd%��Y��?I�Y�U[J�Bt�kr/��HG;�C�����cm���߹"�wιa����&Z�ᔓ�̛֬~*=�x�4*UxҊ������Q�$�a��Y��:�?@+�p��>�W?�fU�я�.�=��2�p���L{�J�#~��K��i�{`s_�;�ۚ*<�όx~ظ�'fq�rW6[l���u�6G��Gm�?�\A|��Y�SLX�
��'b5!�|�H[��-�l��hY�SY��y� ��X�a�0�ը���8��Ba%��b)U�fϙ�'�ߓ~/.���^EV�x�V@�/�
�^w�u����N���뫮���,���^>���Q � @��#�S.U��o�i�c�°�^KB��ު1 ���\w��`X�p~����-w�{����@B�ΪUOm�M{�_
�M��;��sٞH�C�#��0��qY�������\�a[X�<'	,�/��~�����;��=��!1��f1`��җ�d��3�I�D�ôe��p�J��h��^1׎DB5�bHJJ9�laӭtf�
��BZJ-yC1Z�n� �؜ΰ��Ѝ�T��I� ã�?���B<��Wq!�hFZ���O��-���7�l�n�Wy�w2�V�ZV=�xX�����t��l������T�2n�Zm�E@����L/�0����c�3Ꙕ��p�7K����ņu�CgY��MiqqʤV�6��$q�2B����� |F#x��|�.����t5e����
�Lm�W}�#CuYM�=�C<��"�r�`dl4./�åa�XH͈ޔ�5\F\ �� �M
?QØ�@�P�ƅa|��;�y^�2��z����s�����/��'�c��) Taz�CwO�u�d΍%�nI�4�
�Sփv�k�L���o&)?�4������Z���S���:-�M���v�OWGw�<0��ss�ӀQӖ����4/ݼ�+�s�9���~`�_����芧��֖����K�no�<�4�b����Q��r<�h�1��D�G?6[�5*�ٶ��u;O2�>)e��Z�	`��::��M�_砤����@;���Ë��E���/�x��q$��k���4�+c �Q��e �}�O<�.�E�ڊ�Aӿ�=��Pn�R����`G+{����ʺ6̟7� Vs,�?��tǬ8@;�������M�;��I� �"�Í�"O��$�2 (���#�?���?��?�/|����W��/(���-����S��{�.���6<)Z�C����V��k�eo��������'�������2ۢ�j��;j/(+%��E��*tQ�y���z.�����WCw>#�G���X?ߡ0�a�
ݺ��tu϶�J�fx�����5{j����ua�^;�6�gI���%�R���C女p���+��nV)u�q�psX�vSXs�TI����6�n��=b7�?�b�<n��ִR����t���Ȩ�;�n�.��_�o�}�C��N+\$���e�cnˎ�ɄZ'�TQ���(i��0	�t'�P����ڐ%q��*Y��?�i��xF���O	��`t!�d@���.� Ý$Y�_=Ҝ��-�fT�:�֦�����a}X�~]� \�g����x��C��Y��N4 ���MF�F����	�6�
�V�����{-�#���;�7���W�5�����Īա��k���ƀ�����B[�]K�i��s��VD���p�aO��zsX�a��*����[騄����~����ͻ��s�N$ox�����jx �@l����g�"�EEBB���Ԗ����5/یs�_u���������uM��RW��U�P5mi���j�����\��_���Z�v���-�V�%�<1�j�ق�!v�����I�U��9�<]�O�����{�Wx�oSX�iM6�g���U�[I�ݬ�粽�I���Z>�߰1�u�=F):���d�S�eȚ>몃�?�C³�����Ǎ��'J����3kd8����Z��QO;&�Ǟ����k�F����mA�g=�n����j� H�PZ~���t����-h�Xpmi˶�o���� ��w������y}���z���ʯ���Q;{�_�|��&(o�=*��>�ݴ�8��_g��W(��ܠR��\H��/|���^�2��R�c]�$1��0�|�~��������t���/<����xU2~��v[N{�s��
s�.�c�����]w�6�t��;c��5���T��!�w�WZL~Y\�I�{���|�>�Ʀ��G2g��ea>���ub ��e�p�~���VOa��
�ָ}(�W���:5ߞ�(�����J_O�M7�d�1ա����(��� ���O�H� Ҿ���U��J�����i��R�导� ��9�=�г�q�f�!`���A�0���9>u���W_}u�m�Ea�ys��y���f͞V�z2��m�r���|�5����7��^{ì�9���U���o&iB'����������a�����a��9T�����oF��~�j��FTra@��+v��;��U�<h-�do[vv���
w�[U���o����r����zܨ��0~r�?U��ߛ]�z3�f����z�*�J[7��,���
�b���׿��]�O����(~y@ZL��^~��-�=k^\ ������@�ي�2cq���QGt�u��{��U+-<T�3��m���q���Zޘ�%��/~�?����7�����q��W��6���ׄ��+�巈���������fx���;�>������28���w;�Iy[ڲ�ģ{<���jCi�ݼӮ����m�$���y��6��gaTY\
`Ͱ��l;�W!��"�c~����I'�d�Y��	�b�Q�N��������O<eq'|�;��:t�;(b�i����On��y����S��*�^�7+�R���m��fϝg�W^n�����u���LY6i��?��n�:(-'��!]$�����>����f�q �/\`!{�ψ~�c3,0a _�5=`۲}e���L(��̘������@�u�E��8\�`��vBj�S�UΊW;�ݲc2�Y��r�c�D2t-~��`��>I���_���l���MA'9�o|�F��^Q徘z�B����|�*�n8萃��˖[�?�G'<��#�E`4��\�6ܗ�3�B 0s;y5asey�jg�ǒ������X7��?�x6,2���B�=����W�j�\F�O����
�����G\�mi��*��0��ϕ���	[�V����%�����{.F���O�f��Y�[��A�VT��OA�5x.�³4jBA���O�~�к�{�F� �
���Y���Z����O�G{4k��:+{h�����z���xB�X��}��]�5�`-tf�a�q�ש�Q�d
��J�!i�!�Ց���^X��/�� $9������e��V��(`[L�V�}�X�FZ��w~K�@�������	g!�<��/�	���5�暩�����:�*�B*���{�"X`% ���~};P��HH�}�mn{J����3�Z�V���Xv���ζR��Ŏ�ي%tS��
QV�(�T�b�'�ݡLq��ϊ���H�ߏ�C�{�Ï~�#�ü'����J~r�$����c�CF]�і��7��V�e��vU�F_�P��J�⌝�ʟ�݄m�TMNu�g�k�E�Ɓj^,}�9��L>�z�<H� ���FZ����7�).&c	�X�WyAS]�#XQ"Ucb�
y�y����C��Ct���#�+.�;)�c�>����[�o�_�}*Y�R�o���']F���X�ԓRP� ��^��͏J�¼s�k&�jod �����_�����Ð�}��`��<PO~+䞌�����1�כ�(���?.���Qyc��^ײ�6�^:9�܅b�@�(�z�[�j. �[�����e kLx`�f���N-uo(k/5nbK-�$�G�=��A�K��N�Q��{:�f�Ų�EQߓ�>
j½p�[XB��Z�@-�gX���u����MI���/�B��g����D�@��(} �]�V��9
�3���[���;��1���p4t�J6�E��E#��5��(es"d��>q�_#��j_�̜a�R���w�{T�W�͇?�a3�t}8jd���Y]-;���%���]u��M���p��W�(� ��|��A�í�x}(��hpȂm������0�({�Ϛ*�r�?�V�T/2S�FEp(D�b��𚸈��=^�Π��E��<(zAh�e�6F)�d|�����I����ڱ�A�����D�_�GJʟ��$eP��@%>(�8I��WD��͵���ͱO��fVO��V�Ŗ�R�fd�o�3�<7]SY����~�%�Y#�Zy`<��m��fc�^��k�u� MhgFf��yK��rke�+�Z��/^�r�/p��`<��ۥp�&D�%$&?�#�`��R@^���5�e�*l#��lb���>�*�U�Vc��-�֥ב��B�d��R<\JQ������^�F~�����Pl&/y##0�P��țsF�)l%Ũb*?~�@d���K�Y�v���&��l��ª����Q�@�t�t�b��+Ua������Gख़��gˀVV��f4��6���暊��z���sm��3����tq��W����V�~������R����uq6?��=��?�IG�&-����($��m6)E'%���>�z�>�.Z1�k��&G&�X�:�֑Gi
��@��>���}�/�]�\�ue1s��7�Z>���H����
e"�N�FU���0$����jH�Q��������1L��������<\�7m���I+��c�!/Y��pH�o���?��&a;o4H�3��a~�9�;ƒ�����FyzJ��#-*�Qa��s�O2q�~��W�IǺ�z/r~c�(H�,�}�))�)��G!yإ�<gx+�_�c�X0��؄��,�~eD��M�䔬���I�s\�dI�O�gAn��Ip>'�A�)�t=��gk������,�f��ZȔpTX��%�s���t�:�9'�!#�EC��z�#�����M�K?#�~�;JF�2589�]���,5lJY���Y�w���04�.�T��0����tTlQiz�uBz���jg�j���9���t�VR�Q��ku��ʴW���8�}�Qc}�V�����z)g%"�KO�UB���C�DV"x��+7����?
DI-����1��krj�q�b3-R��z�rC��5cA=K�ԑ͔��x:&ŏ9V�[H$��PD
1�D6��;j(�筧�{�~GAWh��=��A#��b]K���Q��(�;�<�&���`S�V�J�S�HcEH1�-���܄�Ac��W3=�~kԱ��fe�Q{���к�J3�߬·R�j8�a��ڪZ�IȔ��:-'O-B�db�zG�k�'��/�������ڷ��5����J $q$pa3��w��h��0)�=��::Owg���j�����5l�^i������2���#-*����^�h�q_�&���r�0���=e�g�CǪ�i���PЊ�9��E��YH�63^�o�;
����N��!;ϸpu���?d�,�t)�Q����@H�{�+]'��3؊95��0VA&Ǖ�sOZxձ/�0�E�;�.�nʍCc
�:�s�OǤ�u4�Oc��i���a�&�c��]w5*VU�z��Q�d78M�=Q�����h&��w���o�a��e��
ӣo�(�&�b�<� դUa����)�YY8R�,��$��ީ�gx,�����'/O�s&�
�
!�R&��QQ�����ߔ���(�z����^�+��<�Ƃ��p��<U�1�h|)�%e��������RE�'#�X��?�C���?olճ�uZ���e�]L���	՟�Z�9�:�����PP�'�Y{�4��	a�Y�������?�䨄>Jm�:ʝ��m7?���OJ��P�E���_V�x�]`�KC(�j۷y �}Κ+� �u)b �� �_~y>0&�:�.�&.�L���g6Pe�kA�v���,]���j�l����W������=TL�
�M�ܟJ�'�T�7�wW3"��b�0c�q�x� Y�Eԙ�c�#)�E~"D	LY���9yT�Dqr���sնx�׻���TG)�V��/��\�Ej�:�K.&x՛�!5M<G
�)�$���+�cW��y�ᤓV�=��==�J�7�m��Px�Ǭ����z�Ø�[XX�ɴW����]mC��3�8I����n����M�q5N3�==i,��U�BϬ��Y0���B~<�I�l 3�T ��&���Am1L\���Kp�f	[m_1��!��������O����b�^� �$��$/�Rca*����(�K�$����Q���E�(�F���R�0�S߂r�a(D! ~ON��2d���z�������﫝sJ�Y��XT���t����W�e1���{x�P��T���q���q$I��!r%[�jIX�d���z�<��p��ׇ+���NW7׫�<i���6��M���I$��N%��o�J]�d
��|����c��@�%�l�ޡo0~?��B�pË��v����D�&�?� Y%*�A��'� ��K���	ca���<|t��欣����u��ӻ�
oy�xkE@�[T� �(j��7����t|��b"EJU�A��X���D�U9	��(��Έ3�3�󂹧0k��TU,�w�qǍ���ʯ+4+��T��74&tnԃ��cn��؇�FOPV�+����ܳ�	'�8!�KI�˥Z��;�d|��q� �6�<�0�<��ʧV�cc[e(�ZCӗ��l	��>��/�ma��w�yG���_��}40�
;����V���?�~'R'7����&�,f�;�!�� 4lrtt�A�i�X"�e�w�.U�
��f�2�����lU�����
1�z
��(>�������M��SY�:&�z�F��>Wa+�����1I�,��_���S&�x!�B�SS�õ������4��&�����3��R��������[��ݏ?.|>��`���o��d�bU��v�iv�4����(s�'�|bڏ ����3���w�֬[�ſ|��ê'�O{�3�ҥ�����-^�]���Ӱnh��e�Z�%cc[�|�֝^�����љ��
+W=���DK�?t�l�bQG�7�p����Uk�QO?6��*�R����N-�<
Y�~Mz�bXF`�{sT���#耱EO�J�AU����G;,|�<����ĳ��8��"R��{x��d�VP�����E���d��ZBQk��W��ZBaފU�x�V�.��'�=m��&�E�|\��Y�F��ys�KKR/�m�������4W��|������}O���Ҽ	����V\��`Q�oi�R����/�{��a]T��w���9,�M}����~���p֙���S�@����([�ʴW��	@1���Ι3;U{�o��M��H�Kw�����?�)~��.�����}���?��!y��7c���z�^hȋO�y6YXF>��cͶ���#4�X4X��,⛅��
p�F�E*O�;ؤ�*\�7��d�Bl���a��yy��M+�UQ�D���J�
�H����"b!-g̞�{�y�Ɵ �����֬��p�C�5��r�~<�Z>^}������o��C�f_��O��p��[N�s�?�lI����
룞Y����_�bx�E�	wYl��#;2<�Уa<-�g���	tW��K���m
s�v�[n�U8���򽉟�5k��;	����as���zVX�nc�����z4�<� m!�x�	<4yx�^`�#{�'�MdYy���������O����C 5Ƚ2���h�d����^���tN�!:��]�"_Q1Vު�ڑ�$�����mC�WJ�U�L3�7�"2�\|ިH���0��[woC�	��d[9~�ܥ�{�dk���И���?�"�EO��^t���1�c98�F�0�U�m֪᷿�9��	a���>4d���ӈ���V�z<>�V>��z�r곭Q�A~�ӛ��F��Z�.ȴW�I#��RͲ�W���3<�أ)�H�ue-�Y��G��ąN�E �o����`g�y���TSx�'���/�5�җ�4��_�e���'ێ�j)�V�r�-,N��aq��M=�d[�SY|�{�e��D��?��Qdx����˛$L���ӱN� y���i�B����~���r�O<�8��
�%��@�+W��{�p��ˣ�9/.��3�� J�[�TaRl�J��<��,���.��#�?��p+���W���PO�B�ء,�����!+��������>��+Z!�ërχ|'�/I,P
,x~G�׿��f	(^���b���M�����+c���V8g\e�QԬF��9��'ק��L�թ��D�PR
��o�C���y
)��~����/.J��0�"O�WI+<Hn���%��+����}���Q�j�ĸ�GT��
�R�3�W:�EtpB�8�fu�����A�E���<�#�^����jQV�j�u��7����՟X�]�ܙ%]C�����qM�:�8�,wA=>a���ĘZ���7B�8U*�jB�4�!w+�˒Ŝ#�gC6�ERS=��E
��'baf,���~�|�m��62
�Qb#�0��&Y���IǦ� ���檼`<\B?��Q���+�'�=x-�a����\\l���e���`^w�Q���OL�uk���W��ು�ƥ����[ݳ���`�YJ%�!�^*u�M*UR^n"�{!atS�^���O��2�L�>�{���y��U�F�8�BGE�f�E���L�\�ĥ3�K^���O~Ұ� '�˼=e�A߶�GDʟP�^O���Cё����~fFA��B񵒱�C@�`
���G�&��	'�`s[ʜE�ӷ�������T�������ƅ�V6�r�_�V`��j�~{��.:�3�#
�&���L�z&}�tRp�kf�ww͊�¡��Fk}m�Y��h�f�QBgX�;�Ǯ�W���?�'}�Ї>d�>&(�?x j�۫ց�(�y*%�&+b4T!�K�[U�;j�E�����F��-*��)  �G90U$���J�W�J�z��b�Ó��]:v��!� ����Kx�0F�(:'e����9�ȧ���k��5���:u�9���u����-�bŊlA������UO�L3���	�j��O��]ʉ�3���{Pxr�C��G�aH��*�P����[������ ���Zgq�f�q��)��(8٧>��N)@�>	5��2��l'%(�O�xK��
�R[;�0QhB2�^�>�-��4��c,����\�\�o��2�h�񊮗�E4J���Q�V�}��P��u��4�p��>���'<��á .��]�E	�gO���ݢ�K�,��E��v0b^H��<M9"�T�_ٴW����#��}�s^�={��5�+,�.�~���~���Ҙyq�8���1ǝ:����V�V���
_��YU	"ڽa񫠊���<jH��2A�Of�_��2�t�bX�8����w�(�;��d�c�|��4变r���ɂ��fAP������@�I�&���������������}����k3 i;��cC�^{Z���ݖ��_���0ؿٸ�6m���ts�qǞ�v�3��p��	�@J��3*�g.�O�2��:+�B��������0{ޢ��!G�E��m�;V\n�.w5���h�@�I%7���d ��ӟ��n�����  ~� Ą(E�KJ����SF䕨���b�0����D������־�4�CV�����lq��
������A�|�q��L���D�w���	>=���¼{e��KϷ@�v���s��>Av��n
#z�~���1��%���·{ "��>!���Q�0>��������]w�i�Ϳ��?��N�,�T�` 1�1��$�İ/`�%M���G��M�
!�k�C�3�f|݊���wb��Sqt�d��zvO�O�����X��w��k�i�j�A%��aNT��.�?�x��E�=w���:��|�!)d��6n�W�ϕ�_c��]��{+3��O����K�f4��=[��Z3����h�����E�ȨU5��j�0�:���M�!\pAx��^��o�&\q��k_��YLLmW1Q�&k�S�>b�����K�"��k&n9^xb�hdbiۂ��կ!��j���I�ce��NQ��s£)�*�@�d#��+�b��c���$�}G�yOD��"+��'���WwM�P�B��E�+��B�B/�h��_�<�����@B8��������E�r�,
R�x�į/�����;�1�c����)��H�D�9�1����s���crO�f��o��`*����d�׊sa?P��M����4��/_ȋQ�󊗽܎o�Ż�9s���?$<s�)mC��>�9�P� І�%���)4�zjB)#�O�z֩,J�:_է�7��$(�!_@�]Y)bGT�NJ�6��`�Il����@r���>` ��\��p�r����0Y�-�˕U�;߃�.J��	Cų��H������{r�RZ:�S�B�Hd=QX��/R�οނQ�.�G�����ENVe=���}�zh��q0V�@*���+�}��Z�@,[�0�}�7�*c���£�������LfOx�P|��zECq�T�KIm�k�����~��_<�@;g#|G�~�Be��wA{H���CW�f�q.ox��E�C,<���/�\�1(P� ��K�~��~z8ꨣ�;Jx~)^3���/䞆�Ȍ%v�����WX��z�M7�
#i<ł��Z!��TYV�D����o?+�Fi��]v�e�\�w���h'E�+\�5�Ӕ2�I�q�9�+_��m˔t�:�!0�Aqބ��;����;L���t0�\�Rǣ�g�{˓�c����(���̹�]����X���z0Cmϓ�),e�C2��T u���gE��!U\ �u(�(�;�qSj-����3�Q��\s���/Xؾ�	�
�"�f������?�+Xy8@�Qp֭���	�O���Y �sl?ߕ{�x�o����g���O�$�'bM�}��,,X�Z��6�	p��싱��x���x򋱮�t��w,:��X���g�5C�Z��`�q=�y��F��Ɍ�zZ�Dq�
kEn�o�"�M��h���{��)��b|>
�N�@�L�`Q��m-��@�M���w�-&���x�O~�܂`���/�{�7V>��$

YҜ��d�� N��eeyŞW �}Ja).�܃����X����+9=�2Tx̋�ڢR��)T��o��d�_�t>~�-��Ň�t>�影Qצ�IP¬�Q��΢ �C]W�	{0�x-CB�E�Oޯ���<y}�7�a#o��Ʊ�m��x��[����2�ѥ������m�$�6ʱ��x ��?����{��^{�:�	�1�(��A�����9�ЖI����3~�G��c�'���C�EI=]\YA
mx������c4W	J���X�X*��b�a��O֤� S[;3�G�_)|3�'��%��%7ٷ{�y��XM����x��5X��GǨ��rqY[���4pM��G�z���U�P�6R�XO�c��ݓ+(�O��ׄ�qY�+�~�H<��,:)1�g���|2��̞~z,eQ�#��Z�-�~z����w��[�K
VcH��C�}���3�SCH��@ʠ�exCL9,>c�1t�����Ka�H}��G�t���9/�/0w��_��WٱC�v����X5�}N�/�X�bDe[\C�O��P�)%��6�><���ذO�q���|#����nAt�"�|q�@#%��.��P��J�MF�Y�?ɋ�d�MB���)��OhY%rk-ќQ:�[ ��z�%�BԾ��P-Z]�da!����?�SM���J����$X9f�l�� ���D0� ��x+�uU��{����Qܗ����a����l�+FΟI�dS�h��'Q�,��(/ΗEoO�J�EPJSR/���ל}���kxl��d趾��ay�׍k�}��5��uQ�����cD6�[J����!$��'�M
�Ѥh�țf�a5��߶��·	������K1yY�7�ٟ���;�7\3§�w>������w�Q��uև�Y�Q�Ωt�s�y7{�\�� �cp6�z��a�&��\`o�!B�ԋ��X�B<�#�G��� D���`>~�d�,���QP�E
PP7<�I>a+/AJD������}�Rg�qFn��!��J�Q���cb`��!�K����-������^JL��(Y�LL��e>���d��Zם�1�u�@��mOׁk&��~�m���|�3��/6����d
�Ca��C�0Iz^{@?�|���X
�#�|e�)<H�k�H8��
s� ���J����'��SO=�ƙ��
E�K��s���k���4�4�=�*���xd�(SZ�8O�����d�)��v�NT��%ijOpj��a�>8G��]�앰ւ�ךk���n@縵R��8�������U6�����2R�>��x���b� �()[M\�A9�*B2%KE�X�P���ؒU?9�ө���R*��� U3���ۿ5�Id�*�^�W���T��hC	̕���Q����(��4[�t<��|�+��ҹj��9�""h2E��#�J�^0J��9�z�ߏMY��������gD^'���'>a'��v�(k�G��vAa�X\r�%f�{�[�iy��7���"��BCR��X�}D<�Ya%b�,:��\�����{!EM��d29��H$�-��_�a'?������Y����Lsр&~��镧���y<dybrJ��5p������Ʊ�� ���#���N����{�]w�n�_ F�m�]n�$��R��`��*(~Vᕼ�}�3dぞ�J�+�Ȃ�� ��N*�=�n���9:�f��q~��"�?�S�I���V:V-��/�5�����%��-�j^���,s�÷��"� ��R�4%�j[v�裏��|��W�DM�g'�t���p�KɃ� D �������*�$i+�F2�y%wQt,v����{����o�KȊW�/��bJ� ϕx4��%����Dj#�6��^"�<���#EĘ�e�����'j��v)��\�;�5�\����CM�Da�Md��Z݊댧���
eP��"IG|]�p��y�"l�U)�c[�7ҙ�������X�BQ���R	b[�����A
�)�%�4��fA:6���Ci�UO��	��|�BB�7�Rj�����
�u�%n694h}�M�6�+��F������*�qP�O�KK�3�U-�_�1S�L��>mIe[c�8v�R%����ڗ{�g(
�~*[A�YӢJy���C@��e��Q6�3l,��k��������ߓ��WS��Nŏ$�����Ҵ7�(V-1H�C��U�XWL\�4)���~�����b�m����ZX�@�����(�w��?�m�Qm��(Y�L���,��s�U�3�����a@���E��1���Çu�:>�x�0�_,����\xα���y����D=T�T�i���{�_� T�3������^n�{_4�s�Ө}���Ry0�<N;�ܪ�ّE���J㷼�-�}�z�8�[��m�6Q�{"�` ����+_�J��!�O|߃�(���/�+����R����B-�����q��m`xlM/�F�P�^��TV�ȴW��=�o�!g�D�z�*��!FK�"b����CDV��T2�Α�,�?������\�h<��x-cS[ƖV8{Z:�H�׼�5�ȧ��<�*h՗ZL�(�������s��/��3Qt��G�ÃT�f�*�Y��yHo#)r yU������/	Q��2�?@'�����d�Ax�5��0�ô�s	���	5�:���B{��G!(�6؟&ߨ������6�,��a���>=����d�����o_�p͵�U�O�tWg�q������MZr ����+?&D�i��&؃���[[W�R����B��b4<h|M~������X2�Ǌ_(���
K�"����`�\��j[������(�ָ}Cx�����k�r�=N��y b�_08Ny�~�C'|~�G��A�!Z T9��=��XX�,>$�	E��R����G���������Sjܔ��Tf��/%;�寄����!zx%!b��Jx�b?ȥT��e���-�&�`z��9���"���B�!o����G����.E1���6a�f���bbX���)���R��<Q��W%F��4O��b&���������o��
ay"E_��{,���C*�!���������X����u�[��Vر�xE�%�N+�B�o�<�?F`؉E�@�T��^
����ʁ+�䘚ë+������9dWPȂb����rDC��[c�f��I��}c�q�>o��V;z��H�n7�0��m$�ے���3x. H��o�h�IE�+���}�E�����ٶZ�"���V�%�g�D���E��_�%j\� 
���k^͇<���rQ����+�s�8�����M\vV�ǟ���ʿh��l7Ӈh'[!,!^snX_|���'�{<N�X���˲?��g���|vu�\G�F�o�zƭSA�=�xA6Fs��E���7��DSma�;�!h&r�Ց�S;p}��s�?�g[R�u��1(G�X��ͮ� �,�,�(Y�� �4��<+�((*�����18 ��,�Z %�C~�Lh��&d�3���2ɇ)?��T���(�ڷ���ۙ%���TM{��lugV���n�s)��9_Q�X'
Z�Lաk�I
���iʚm͝=ǬtQ8�j:=�����r�-��ũ�dR<ZU���X�g�u�uR"�� ~x��!�Z�#+�,Ă*ب�rK�E`��/Xo�Ḋ���U�3ް�?��O�7�����_��_�؅�����YX�4Ua|���4�-�U^$h1�Gq4)���2��1I:�!��7F�ƫX8U�"�-Q��z�m≰�����_)猻;��k�TJ����������Q|��^���M_��}�K�o\V\]�$s�`�z��>���d��
b)
��@Lo��f��O,�F�����!V��a7�/y[=g�IQ�y=�>��R�x��IֻN��#Dm�X��(.:tѪ%���7�$���XM�W�1n̂��@�?1��lC�Xǀ�[�2�+'����u��	H&���DH�?IGwG��ŴW�q�k��������I%����'��-Z�>���dՖ��N%ٔ�U��1}�6D��Ќ�5�W��U�Țc1�dl$�0<��9�Q��W�V�~݄�����L�o$j��ppO�N�?��8��҇�9�I��C��#���F�TM�Xt�z̿��=�� lKy.O�k�&C�J�<Ť�3��.�b�?�fo�K�B.�X�r�5i4@}`O���C���)���7�֢��M����ĵ���\CV�g�(�3AU��X�R^����D�阽���,E˾���S�Һb2k��ux�8�h���W�D�"P�9�43 CUOy �k�Lݷ<�ƷBA2<|����YO���VD��+#�-wf�T��==s���ٴW��Ty�[�^	*�3�E3$#�gE.M�9����D�)�llk�%!�����xeQ��E֥�s��e�Y~!Cl���6��˛%�&�/
�
����+<!k��J����\C*TI(*	�1#��S��s~?���י�&	UOR���:��"f�b=�>�\�:O�_a��G��O+���U;Ey�y&zD����n ���$��Z��K#�?U��E4n��"���_{?G4�$;��/gƛBV�����{.YR� �ښod�����7͟?��M�Ԓdf��+��H�Q���׾6\t�E�$D��r~��sP <�LEbp���z��$�'��T����b"���7��h9u@Sӟ��!�g�#��8F���Y��9%�E�,�&�4�t}�U�:MT��<:mp�����\�׽�u6>�؅n^���ã�?6�8i�։<o�5����ق�n�=������O��{�d�ƍ��w�&�T���D�&%���Lpoa1�9a���Ț���@�(!rI��	���g��_�z����R)ԉTVń�Be`�9,y.$79~�!�bƱ�:Y!���3Q�L�+��W��ն/q�����h� ����7j���˾�e�m�ehK#Q"]p�Y�O~��+��v�+���-��Z�7^�C�"k˶��1`���y�ؼ����b��C��v)U�i17�p���k� CNm�JHM,A'�'�^��c�'�������
˱ `q�|W��^��(�a����J"��K/5���������}�5�� ��7����>6�����!�EcY9�ٳf�{��'�-Ӟ�����O��v�i���\��5ض�'f[FD�F5�'!t��=R�R������ʿ��  �IDATK|<_}x��Ǫ�E����C$F[BO�ࡒ%EZc�&�΢0�^Z�|�J�m�d	��ZQ��9��0|��9F��.��2k���9v ���+̪�C߄�[{N�.�gK�-���u�p��ϸ�W}��o���GN?���]u��/]�p��(+� �k˶��v�!t���A��4)N�EL��_Oi��P%�s�,F*�����{,dB�����o�=��_,�B�������*����.�U���eL	j) <�n\S��e�b�E��G޺�0��x[K���CG<�w���������W+N:��xa�V����.�BJ8*$E]J�����x$�^���#Z8>
�(tCD1�r����%�&%E̽M%��P�6���
�����VHj,%:Q��J|q�GSi��?���jKt���el�H7�`�{/[��?��?�g����~��߽�_?;��T�����˷'[�dbЩ��j�	��LLe�'��)&�z�h�Dr��5�����)�9L�xxa���'^W��ؿ�f��F�Χ�5�����ب�=��S�s�i��q�����ZX5�5DiKs��F�E���U�|�W�n�(�s^�������>��p��܍��L�3�҇z���r���1�})
D� ̻�cҲ�FB#F���g�T�����"��p���#<�J�[����2�$�
u���CY�r�J�������dm�߱@;}���>8g!l��6������p.)�^�~_�s@	�j����}{�"�Aq�~#�c��)�(rA0��]�a}8��s�Yg��~[.��,�_����}g	ܡ�P��W�@��ZĔ+R�]�FW�.uƶƱ�PZ���:-ORM��S�ҟ�\������ ����贿��~�zvϬ[�;�[�v�(���E�\x�_������y!����3n���������Y)�XNr�Q�ziԓC���'V>�+ioU�m�(�,w~���z֞��K!�G0V�/v��C\K���?��k���J��x�a��^���:�!X���ndyRؾ�I!�祰�/L���J��gG������Gы�Mֺ�N�C��Їrg%�=lјѽd~�}������^DcQ�V
�=�P�M��>����<~�,�>G��Fk�#�2e�{ Bu��2��5����.�����6� 9�S���{^o�y�Oc��^��d��j5�h��"��ui��a`���:�+�f��"~�_�x /�1���+W�H1�>Q�)7�S�� �}ݚ����Ś���G�Ņ�,��x��\��r�0-
Z@����/�rjF�_�=�_�I��2�����A�؁x-z_:N]#]��H����s?���=#&"h,�џA���C��gh|	��חmiAW1"�)�HV�Կރ��G��M7ݔ�85o���}��;�h�^1��8���/~�w>��4�݌R�тz��o~�7�x�aq@h�0=��Y1�~D�O�q���R��)��&�,:Y>�z�]�c*���v�R�2(�B2J&2�e]�-��yJB��Q�C�аV=V˵�-�~~�P���Y�=�s`�{�+^a�y0�:�΅B4�g�������0��̈́��,jfy��q�������*�H�PD4��Aޙ@��}���c�,7VaZh�D�x�Ɍ�Y���&|}�T塘�5���C��3�<���og��G.���?��ˢ����'Ƈo�T�鞙����Wq�vu��1֎�&U��\<�rɬ�v��L�<=l��ΏG��~���&�b�b5�����6����{�"�_�I�&��5���-=����
���h��G<��o�鷃�Z������J$��B4�Z0u���4v���Tϓ.BZ=��b�ڎ?�/�k�,�d���l�"_F�����4ߢ�A{�0٩*Zp�O�Hظ�{|����[��S�q���?�㣟�������%Qyv�϶�?O� �#7��S��DO���\T�|�Ᏺ��p��h��Q���G��w�����xp��U�+�h�vw��C��Z-�,�Ks�RZ�aÆ���^��D��v*�k%���TW0^��r�|}��DI���¥~(~y���=%c=ݶ����B.�7n���v�/Nd%�Y���Z.��̍����0v ��xF_��+dO��Yq�Iy�B4iq��i�>�����@Ź,c�'�=/�S]��ո@��q���.�<��ȌS���_���~������V�`�EG�B��ʯ��OZjB�
�sd��z���'�����)��p���|�q�-#):�����̙��W��e�~����c��c)'=IG)�UX����k�w*)���&�Ox*<!�89!!W`�$�O')�<�W�zo�����!�c�9��9�~�Y�
�(ɫs�sy ���/��/_~�G?��w�m���<^��ZT��4 ���X��.��ҷ$õ?�;{�"����:�dF�g-zr�XK}�L�^cYqx�'�����1���Nr�_����h�X1�1�O,�����/|w��[��T���_�����߿��7\s��M�o�T��RXr�YU��M$}֊����2�a�714�O<?�(������q=��������o�г���Uc���]PH�k��{�`m�+$,W�IAR�bŊ�ɷ��,h%=�7�=ďC�p������V�C笐�^�|��7��y�I'���&��骫�z�%�\�!n�q���1d^h�����},_�(�䓻S�D����g��[^��x����/�QP`-�B�y0����P�ђ|���{sl�og��G����7��w�m��6�n:;��]
�zqmo����+�O) ?�䎓��i�mb,��b�԰�jõQ
�Oબ�q��5�dg�GY�x�_�����G�R��0~/#������>��Ǉzd�J���RH�ڄ��zƆ���?��?�Qu�x��Op���;��7\{������x^�c���șI�
e�=���O����ւVTƾ���-��Iw�������]-J��9}�y{���j���6Z��L�D�B���*����y�����[�����~�����-oy�O��M��^T��R����
�Qp�V���sl�뮻.�p��H{����I��W��"���o�#��څ�כ����x�O4���81���>�+���L��^#����Tq��vi��9�3�_y啗���kg<����4+U��\A�+��зU<�����pǈ�{�ޒ�I�W3Δ��h�f�;�!��� FyGq����֊�W\������n˾g��G�K�ȥ��M���OƋ��Ύ��!�Rф:T���PK�\&Kd�kr0@�!x���p�
	��Ysf��j��;n��N�O�&Չ�+tuu�[�[���w�p�	<�y��{��8P�[a�}��YR��r���a���	����7��E[s,�{���/������*q��׻��X�2�a�l�h;��*�v����z��oG����9.���줮'��kL����d��'-��������u�kf �)m�ɛ_��W\q�;���/���G~�O��d~��#'d)7��<���x|AS�2�
u�}&.5��"��Xg���)/�XY'��/���:�c�)~N��؞����}r\q�f��tW�^+�-Z��YO|wQj�$�?��u�\s�����q^����W�σ�+���(K��m(�������#$R����d��z��>
�f������M�q�^�]y�Ag���l+'�w�����y�{����\saT!�tw/����Cx�f�{{����ng�q�s�����y��Y�U1�r#�6�Y4;�fʩ�ҁ%�v�����+_�J�c���8;�.��{�0fY��9�����<�Fֲ���!ت��n�������:{������+�,����#������^�|���H!-e$��x�\&���*e�|R�I����h�<�`���8a�G��w����}n��n+�:��������ݯy�k�sϽ��q(ύ7�8��;Z�'���|��P��^\����M����m�������ۗ/����u�Y���ٽ��.�&�&s��=��me��]<��O?�l�n���mrmN?��M�������O��O�|����&"i�p���P:R���h㦈������1�&������=��1������ӎ���ۿ���+���}�����?+ޭ�{�����7���#������{��7g�x�:';��	�T��	���|�é%�QU�B�H�5I��3�C#�+_��׿+Z�+C��z��Z�kD����+��s)�����a!FY�8�c��ړa,�����>���;����x��ZI��"���7�a��o=����-�&W4�8&<�x�6Ɨ���g�]��O������{����	�w[�� o{���>���~��{�%��y�Q����dxy\v���0]���WI$CV~R*���L.8����YSa��JI�aҷysR��`F��,,g�rV
S.�=���R*ل��;R�YRuk�4�`pB��RP��;E%b�����y�m���@���x�?�;g�G�F�#��wߓO<��/�.]J�w��Y�f͉(�6'������q(��bի�#Wz���z��Fp�Xyka��%�F����x��h�sSk���^o�F�go����9ȧz�Wuu^�ˮq��R�G�X;���@�}��J�8G������m'ʽUʕ�;*b���Qf����8�x惵�����rg�(���R�RI�zŗꎇ�}����'�\J[ܛ�{T����j_<��{�������C:�8����7��(m�������W]uUwTB��гf͚Yq0΍�DԡS8�y\��%j%dcJ�n��f+��w������7�3N�2Ǥ��5Ǥ��/����&�4��1��uR��'������~v,���qL|���K�������x�~W�Egէ>���ƒ�x≏���?�hT������R��n^�#�e�m��3>*<w�7�d��g�W��H���Low<^����.���,����w	r]�d�Prz�K��^Jo���&��4����@��@�����uB3�;�Z�T��{���;z�I��ܶ�1�W�XfPƱ�~�u����gOs�1�V.��~z�;����y��ٳg/�ے���.u-;^�A5~n��{:���������k6��㸩e�|>_�h��yvM�l��`���K�=*�����54��M�D�%��&��9r<�cw .��K�,�׭wٲek�9���7�%m�?9�l˶�
m��r�i�Q�{O�d�&�(o*������k��Z�%�z׻n�nm٩����ҖqH�M�J�������[�Җ��@i+����-m���V�miK[�2����Җ��eJ[���-mi����oK[�Җ(m�ߖ���-3P�ʿ-miK[f����^��2�R    IEND�B`�PK   ���Xwt]i�3  �7  /   images/612d2f36-6902-467f-9552-2a5db1e13335.png�{gT�[�n@��(�!�^��Q��ń^�Ы���@�*�"%B�UD�@�(5T�����w�=���c\�Y��s��������}��Bv��"SSU���� ���+@��c��뺛��D�N����2� FjP5�G�k�	�!�%�">tD���e��?ie�cI�'��������_ߗ@����
ts韴8�/"�*�H���򉞂��g���xع��7ܪz�n3�Ҕ�qu�~�����������$�t����|��\<$}dX�Ԑ҄l>�?U`�2,FZO�\�!L�����,�7�����_B%u��i<ɰ��`n�||��޼�B���||��|��`����f�v�`������q�w�ٻ�0��_�z�dXX������A|��=���?b�J�x����oB��\ɧ�>'cE{g@=��B��|�c��������������R�����d��2�4�υ�R����������eoH��ǚ�ި����PS|��'k}��Ϛ�-�k����o��]{C�m�LA��-U����[�>����b�3����QW��>�1�âw!�Lk�	 "6�D;�)�u��S���++�K�{������VI.�����1���`C��C�A���+m��k��]�i���/�����2�%�_j� S��M
UQU}s�KW1���ғ���Ы��H?_9�N����mTTR���O��+h����jG����������|(0�K�%A�r3�[E����#I�}����|��QJZZ./H�U�=�ø��[��^���n��{�ﻳH{�tv����\�[�}�y�{�~��t��q��f��FM]��c�QC���6����U����N�N�$�?|�,c���2~���&�p�Q���m�t{&z�*L���ݚ<����� OOO'�nwD���l�Z$^�� �#$Jb�JO���,?c�phe��*��{i����!�ߨ�����-s�V�|9�G۽|�A ����I�R؏6������ZI��z�t�Q��`��	���{J�8T�L�܎�>Fh�R�4Xw�������h�S�/�0-7��NJ��A)��n�[�����D�q��]�����F��:�U�<��2���·����m̏Uk����ڲ�}&l'��]a��\��`ڟ��EH�Y�#F�f9~x��666U�Ġ���j(	B:�x���o�璠c���k]��$�mW�0���.�gǺ
k�bo�U���l�L!��c���c��+�Yz�wy�ֻ#a+��vl9������>	� �,��,m�3�=Q��h(���A	k�u�f���پ��E��g�D�l���d��4x�b��׆��|-�bh��KN-91k�y��3Kt�+�/Ƹ��Ǔ�X��W�l��=�	\9���;Z6�.�]��ݜ�>��S�C�j���9�cئ�K��B\��zjg��X�	6�ᒒ�?Z'wq�S�:#��F��D'�z3�Pa������zc�O����@ +�x��7��g�����=�����=��_m�MS��<� 9zr��*���}�)`{]���O�(;�m�O}~�Ղs� ���m��<jZ@��S�7�=�~�Wd�NjS�_Es�܋���&}Ox�k�e&Ղ7�W��uu⽛X�����O84�4K&V�JĪ�\Fj�����*��r9���������p���et���B��((��Q��g)7����'I��pG�e�䶇�M�	�᪻ұv���@�b�د��X�V�c�A�s2�V��KWM�m��<WRb�	�7�'=3�#�V�_C#P���tĕ���ބ�����
L�>m�Z ��&� �qv N@/��
�=y�>Q���u*�`�)��ق ��U�;��C�~D�K'괼%Y�活<�˪1���J�*�>Y�Q��>��_�dPIQ �zh�[R�M��	������r^�IC�"AIE5�j#����,pLA�/��f,YG1�j��g�#I\G"4��~�ȪМǟ�x^8��^�����}|Z�@�}�za�0򑀛m 8t�qx�+(,���c��r���Ӎ�M{ �� ���Qa�p!1X
�Je���5|?��ay¤�3��%4��KIX4:O��U�';�b��C�
s��.فoUO�W�M�CՅ��4��M��+�z]@��O�\���i�7GD�Z##�ks���ls�h��ڧj:Vn��r Gp
��G�mN���pƢ��F��U��F� �Y���﭂e�
o����H�+H�<�h�r�O{�j���K�A E
��S7E����&������� �.�B�����EFZ�ْ����^�T �J`�RzB��YvW<�C�mD���Y��X�z��M�'"���9�g&��C |�nu�ޜ�+��.
rk:*@�Bz�7��Z���3��A���5R̰XW��7b�"F۶�5|�@w�7���5�x��<��ҁ���J\�W�B�ML2�bب��1uFN�>����@�����<��m��l$���@���3D�6�r
�6���ɔ����&Є���&nmk�ν��u�8�(o�,$[X9�Hʁs�f����T팸�̢p�`k
��]-���tNy��2�.Qq�'Q�~����\�А��]��4���3k�{nw��aF���6�s�&�7��-�����e���8R�= O9�𙘼��
���`]�Ճ|�^�JJOX\\�Y?����[a��4aaaaKLG~-O�D�9�z.�݈O�b�M�z�En���͡�<�!������2��]M]}�Ǚ��"om���
<��l넶��7�IH�6 �_�ɿ���)_���� <��w#��ky0X0 �m��U���M�o߾M�ΖT��I��謹��[�}A��� �ӛ�A6�)E���&�����f�7��T;��
�K��]���ܬs6�^�{,�U;Ҋ�d[+;ƒ~�t�?v>��d1]{��uʖy"�(v�H�G؞7Dn���h�����f󁺓S���5l�N�|���k���@1�?�}��P�� ��F0���8^�s�ZJ.]E<�Ҭ�oda����?��s�խ�{V�Z��&(8toA�����v��5 Y��|�r�����z���Lm����ŚB�F7�\�[2��檽�t�r���=t����93SW���R��{hZe���-9����,h�w�<ǥ�kgl��)�Ԋ�x���`>�,ll�-��ܘ}�P�Y�׷�����+�7�_�٘j��6Y���ɺ���u�nKt�������b�<��j�՞�ٰ�<]aJ�]@z�7��8Vj����7=�6Z	����KMk7"p�ƀ}����k�&*�SV�	j��v��*�����f���-�Ok��k�p�w���U��~�,|��s�jz�S�S*�� �yN|����x����*mc/Ɏ"V��ub�m; /��l�t\A_���;Ûʖu^��ܿ9���:H��C<����Iz}����x�]�ΘD�"N�Y�f�.q:�tX4�1�c@ȤZ]Q0�C�P�k಴�u=�Km<i�/Z��&U?�>��nD��Y�^�SŽo�Cc��8�g�`d�zqV^G��|��2�I��Q�=����R��}��@U��R%;�Hh@@�����yK~1e�)Yj�B�����u�b�{3n�471pXS���a+ZV�E.�]!Q��8$s
24ȈN��~����Nlz���[5[ғM �������QQ�ס�\����gP"��S��}ֶ�8�a�i��f陥��d֖�!����/�!�K����zG��@��T׶��Sm"��¦�
�$>�
��u�����I �i��PS�:��˱�7&�o����L�b�^�j���4fa�3Ρ�7��E��ts�`m�x�Īu�w8)�'[�G��6c��$j�ۯ䥄�zA-�ݕZ��M5�� ZK�-1�J�b�͍<�cU�K!�t�g���(���CًSԆ^��~7x�u�� zT���n�%O�Uή}�T�R��^|S�IC�����r��iM���bݖ�)�$�"�8A���58��l_��=N%���V��ƱtVB�2�x�֍��^��f�:��"�ƫ�;�d� ��ƴ�����q�6��U��Jy`j�Ꚛ1����ޣ%�|���1����f��\y#boL�E�U�Q^����%<F�f#v$� őB��{�����5cw
d�z�ڿ��̓ c!u;����%}l��.`����@$�Eu�f�_���68S����DMY��d�X�
��
���,�^��)�\�.�k�~V�y\ړ�MEx��9xe��]����<�\Yw�������{��P5�cǭk�=�X[q�`¼f�XS>�-C��BUw"�-WT�
��LD�e��&0+���%\���w'��n�D��������'�S�?�lN��@�-���������'j���\Jet-M<�Y��^��~��39��񡘲Pc��M`����d�$,�0>���������3]=�X�F0e�*�.i)�,�6���&Jf���"]��oS0!�ˀ�! ��ol�A[�;�̔>�� $��ߥ?�ӟYQ���z��j��/~A������4�2��Ϸ�gaWXX� u��"Q��.��V�C>
�e��8��YROF���}=����b����谙�s7�b�YT�\��a9~u�^�9)Ԁǭ���\4�ɲ�fIr�2�$YƳ��{;N�ZS[�d��KrS�'5o̘M�U+�p���qbZ0�J|C��S�	�K\�?�[�� * ]��2��j4Ӝ{�ד��wU(	��k�����R�ҿ��a�[��-��*m�^,�5++q�!/AS����������8��t�;�׫�\��P����+�2�XPp|�IS��R�a���0RK�������&(oj���v���H{�5���M�K�-&�R�>�A��J &�ۘO�'D�i*�(.Y^b@�y�v+����eR�Kk,I^��Bt#bW!8�y���[b?��<�����!������1^��@�ݾ˥���s��~�DmW͓��V6P������"5݊u��qo�i���N[{�c��rF �{�	��^В{'�����+5�Z
'�ʐJk^j�N-kt[r�\�i��lw�&��\Z��&�S�Q�0	����0��+xt=A!y&1�J�d>�={�|�F�}~��v�}���I�ũ����x�St���%=p��Na�QzTK}�^K��OueN�v�:|�ٚ~��a���7�y����.B_���d�hJ*�ނ�{�/�K6�/���Q���o�c�מ�wx�d
�lɦ3^���B�7�B��q�ʂ�L˕+J��l�\卩%W�`��G��[4�4�[�6}I�����^{:�6�<Ș~*L8�?jͧ%�|�2�.���^�R�d�v��sw�լ6�z��=o�b����/;��M{G�Z���l���θ��_�}�@�,�wA�!�;����`�~��a�h��'Ø�!J��|����B;"��EM���=v�����Ю�l ��33T~���Xy���|v�&m�ϔY�A�3�W��2<�+�>�$�Of(��'�Q�t:�)6�S�|�'��8O�u�8_����p�\���}�i����nH{`�ePV�|��oa/�
�*�.&cy+�2�C�ך}��+k:�1��y�E��R����F��k5nt���4��rʴ�o�X����J����Z69G��3����	��)i��O6��>�^���^�f�tں3��#gd��x�~F&c���X<����1[��(\c����P�53�K�Z�m�X�6ȍ%�X�{q�Gs�F�=�x��呁�"u� kƜ�|/���`��l��L�KJ!^�!��|�-��;��.ckO��,�d����c}��(��h݊	ֈ�d��ʙ�XS��F�\M�ka�`JS��F�,���,d��7o�*<6۴���%I^)a�������o�'q�6&����uE�#��S4`����p���y���}��\>���_r�f�H�������`��:m�9�9V����X� r�Z���p�}ۣ��6�6�,Z����Z2��X_�o'J��s3�N�S����Z��@�p>@��y���#l���,�Y��?�ڋ���݆	o,:�hY�E���.h�m��*�g���>�W��@;����Ԣ��zƆ��|��Ӑ���l�e���<�L�/��?�]��:�p�C6�x���R���_A}4?Io�@N;N�����\�FZ�o���N�jx��PD�׶)�g�������Y�������U�xx9���)��4�H��sv�#�N�����2��Uԙ�Z�Y�oHO��9�z2��~	3hV�D�ꠤ�J����3%�ě^O��s�|nHe����
/���s��R\Ξ8JNqp+įV_�^H��?U�E1 �Z*���4^��eF�<33��Z�E�ss��G_k �H������z�5����~	�z�a���qt��@�n�^wOWl�v6�sV� SG,b��5�\�k�8�>c�Z%:SRqʛ��K�����8Y�[� 为D�°ZcSZ,�_[�6ƬK��YG�e���N0uW_�����0Ċ�EV�բ=�^�4�g4�}�l��bڶ�]�v�Zw��K8���5\�5�8MP�u`$�ٗo��M�//�^E�EjX�����;0?�&���n��_:���Vpc��
c�yu��[�e�u���hF3|t]+̸�Ѵ�yf��i�)1�w��"S��q� ]�Txs�G��6x�>P˟�8��q�'�iXv��)��u�ǀ�����j>�m[�������+]R�	te9���bpB{ �߮���.P�^����(ֆ��Ր��j>���11?��8 f����}��:��P����<T��7�����]|֌�0B���\1��
p��X{�q{pw3�N8 �U������v7 8�V�~V`ԫ�UЀv�)�;�����CHf�����y��)�dUc�?���/W�y>,���{ؗ�mu�F_� �(�f2��8�O��H��#���0E�kNU��u�$�d�ֽ�R�G��̽�?B�D�5%2+��!;?kyvy:y����C:e�+Vh&x�FI�8��(�W8�[16?�3��0s��{���,]��ý*#�ݢ��"��r^�_U"^��Kn�8_�?����}�8�iO�3{��	�`)�q�]{5���-萱���^�l�[ r�.c�:��zڃ���P���҈�B�e����)�)�Qpc{���⤣��J�˦^��?j5N��ef�bIǮ߰�5�%Y�߁���r�C�V���tK_@�pUW��}֬�Щ��� I��:6�C�/�~ׅ�Q��9R����V��Bp���P�9�!�])�cX�0�,�m��Ѿk	�]GѼ�!J[�d+�";����tLP<拿]���K�y@�7)u"��¦.��C{\��]�鶧㤃��褌�Ef���@��� n���ϝ(�3�:z�AU��W6����?�O�VzQv�XA���o�ҫ�y`]e7^��>������-|�ˋ�1h%X�+�Ԣ�20���i�"n��I�W�~�eޑͮj{z��c7�t�,Qf��B�'Aq�����B&Lcc��z��ӯ$P�O���v\̈́]��V}��К�j��'[�\�t�5���z�y`zaa��Q�T)l��b�k�Q�A�v~�O�����'"J�*��Ds��{�ϴv�\6����Z�肏�r�
��pfH�T�Fk�onR�,vM�"t�\�p�`_u+�g���ԸoЁ�� AR�Y��_�I��7j{��.
x�PX��ȟk�1���8ß�����^���Ono��3˛xә�C�hM1���*g��/|��;��"�+��p��C��u�\8Z�����o�0DP�H�,�[Y���F`'�.:�S;�u�����#�i=�p�T0��f�ǫ
K�\��VFfkz��hȍ.Ѿl��Q�y'GJ�BJ�+�m���e�G��8�~`S- g��;�&��(��y�T �r��u�K��%#X���b`��T�(�H��WX��)	(P���7��H~ao\:Q�������g��#_Ӕ;�L�w��+(5�Ŧ�i6�+^�Mtm�6-^VV��t��l5��0��gp��œ?jQ��ޯt�
bDȠt�=�{օ��W	�J���u8N���]����b�4���վn�(�
Xh���3��.DF��N�&I蓁��I 8��Tq�l�[9JN�lU���/����Q����#,�����0ْ��P�e�y�e���p�S?������!=p��qwÕ��BnʳW����%Tc��4.�yQRK7�?��Y�b�/��2�JC�q)">�I���*95d+���q:�S.���U1�b�>9S>9�\�f7w�ӟ������@s���RR���63,����wK��6��nH��$]Ѱs�<܍|h��{���64a���x㫜P�c���'v�} b�2x��}>��YB/B��e߀-��8u|<<~)d�/�_0C�<�9�H����� ����D鉗��;ʂش�O�V���{��4
�N�rL�L�2z�H8����[����]~{�dw�[���f���b�maU?I�#jb��qPxŞ�b䖬&��K|M0��#�*Npt��4[��������N������+Ƶ��O��ƴ?:ߒ;�qv����?h�~��5�k ���a)��p�m�-yxϵd1�[Itk^����k�[�~��Q�&]x�(6K��wFj�X��x���ſ�m�9�d���5���5���m�Z"ҩz��s�{t�
0���m=v��s�%�⯪H��&�g��b��[*��cRj���/�*-V�Fb����s,�-@	�%�Yhȿj|tg���`RY
�#1����cg�ޚ�[�at����n��D�ck�k�$hb�>-��f��m�p��dQ5~W�o�����y ��,��N��$N�f��V6�����+�e�\�|Z�[�S�G�Y,��F�p��v��VKh�\�;%~n&���W��Nɳ�=�;'��������_w�[wO"7EE�ˡ����)w�Pl�����N9Ūͅ�|rBǞ��kP �e���H������8��WG�j��@uO�/%��f�������]�(+8/!��ׂ������M����PffJJ�GxC�Ic�i潐���m:���Z�oW'�]�kn���W����]DdDܰf_l�ܠ������	:���(�
bj׺�Mz[s�Ԙugi m�7MCW7�c��bIXg���F��u�#j�Ύ��	(t�Od���pc�<�xx,��IP��Z{l���b;����
[�L����%�z�b��O��o�?w'%'C��+�~~��R�d�ԟ�tĕ�L�_''�)쭵28�+ u��Xn%q{���@r �3A^l���l;�Y�O�@{�e7��a
^�(j�#�)�4Eee��wc<�}��D"Zt�,&j�![�:�r�1�2�̺�G.��8*$�}�_�'O�K�)3�N:?;�������KG!��.��"��#%�R^�<�������I�Ň.��+�"��#DUŔ��Ky��VG��N�V��_a��#�術RR���}���<�a���Ժ�3�ObK��!��_�)t[ RDY��������e�oB�,��ж:Ƶ.Sd(<:��Cʬ[F ��y���؎z���At.�H����!!�g�^�[�; ��x��e?L!dT�c�@i�O��)��u����=�������pP2����������Șf�:��p�}.��ik[��ur9�u#L���xU�BS9Wo�.R�%`ө�(�"���a_'��Q�/��T<Z���-f��G��j�Z�B2���7�¥gV �'t������쿸wu�����.��F~k�-1�*��J������\kì	�T�BMp<Ǳ�+�7��@q_7~�3�7�}�
�οl�F�������k�p)XI�~�!ckk����Y��[O���,;~�жa��g~�L+7�>ܢ⌊���Zx�,�bv���V���D���ڍw_�����CG���g
���1����ǯ_�<ơ�3>|0E��^~���.��%��\E/�|�+i��SdP�u�oO�h�����aO��E���H�۲����?8��xY.�\����%��S��޽K�q`�J��}�Ky�%��}����<��pp�F�;/;��i�-�^l�'�L{5�
�vS-Kd��U�e˾��kqV�L�z����X����Z��
��R"g�j.�����/5��?�ĕ[p�#��UA�Uo�ݽ��k� S[{$)9�0	�
��uL��BT��z-\V�]�'���'�
�cu��g����u�<�خ3�	��&A��*��HMzq���7NI=�X}f�y��#3(h���Z�k/��B
>L�.�u�����\��D��w;}�V��k��� "�
��:b�=�%�VTTzo��F�%<��zOoj����@΃X=��j��ڗ�]���".����-t����[�?��� g��u�g6�l4�5��h^�x�7�7�-���{R�w�(Ӝ�6�=�s9v�	D�3l��y�W�eR�I7�B�jGN��@�^".���P�a[��a5��s�~9Y�J�8&??�����xUq�P窈��W��=�m����S&3�ޗ.`Q�<1� �=�6�Y�W|q�YU؈�ʮN��W6�И#�`�'��-�e1�XC"e��=ш�<�2��b���>�1��l�a���9�6zQJh�և[)���h"�|�IX$�nN�T"�?�<V�L1W8�BDחp�@w�e�cO�d �.a��)�X�8O�`�Jog,���2�v����!���MJ�ܯ���8��כ��-ՁP�p�#�hs�^C��e��dsqdT||Z]����f����93�鷷B���^1_��#)�~�����#(�=333�WSG�Ȝ�8����P�Y��TMLL�\[�}t��h��(�pB��������*|ޔ�m��_�!=F7��:����?J���V)j�;0�71Nvv�f�=B׆=�R^��@��D�4V��M�l��?�T��<ܬ�#E�ڇ26�����h!@ˠ��\�u��&�DS=��s�j����X�����R�1�]!:��v$$Ɔ�Ǆ~�u\�8�VU		���	�����sb�~��)��8͍��Y���}�/y�9��^f��Z�}-uj�j�)B.8(N̸�U� 
5�Z��`S(ޤ�b̜ZfZ[����3���a8����
�U���
�w4�{ǉeHy��a��}��(KKVV��H����'�U�0��wh���lzF=f�6F�k����A+xʭ'�K��G�<��N[� z1dm��W'�N�+O�ﻊ[!���A�ջ���hgK�SqjW��	�� O(@�C�K�|�Ӹ7�:a)�b�>
��H��$�\ı~���¥Ѧ���Pkpp�c:�1�$l9!�N�g�XrBXw-�����Ko��K0p�WE�6�Y���;�J��ƺ��]1��b��������s����愣p1o���d �	�Qr�󣥅��Bz��5:�K��f�/{��F�\E=�ma����?O����В�:2��C�p�=�lI�a{�0`L��_kf��m�e�Ӂ���X-�A1�����靘A��i�ͻ�МQ��������{���Ի�a�:��=\l�m���ar�F�c�q�bہ�ftJav�q�"�����tˠ#$������/\�E����j�-�6����HK�?��ۻ�U��P��Z�����]<���:i,����HGa�5^��իW𙼑G�
����QQ��D>�O���e��c���ʮ�@��?�b�5�bbvWdࡈ!�j����lqY�#�������`S !ہ��Z�Κ�r�
8trx���][�:��wI�
&Թ����á4�^�І������6M����V�򡆛X]:�_�A�>\��������;��\��K���p\[�r,���4�ߙ5��K(�Q��&�A'�~���NN�d(3������%[�z��'�^_�X!�����u`��2�0��S���8��i�-I6V��ݏ̾��*�: ǚY�r@i&�XkY-	��q�D���X ����W��8���E��["#��ǫ{w���Q�ev��� U,t�C��~�7�:R��g�ՄXALD;K�Y�Y}����.2.�%�X�����$�ƴ����ZW��m2[?���0eS�2�/�2g��,WK��a�|�/l���{K��c0���)�g���a=ZV����W�X��4�,��2(3��G7��A�w� �Ǚ[j�z�m�oHx���mMC�Y��V�ioG����d�Pl��Iԭ�ҫw_`�������h%��x����g%�#Mn��������,66B�k��ᶯ��e���-c���Uj��;%�"e�]����}��N���H:���3ؤ*����	��5^��Z~Ps��=�Ĥ���mЕ�����
��5c@C��o��,�ͯܺ��7�c
f��+7_H5��� �5��=�����qd�MO�/#X�=�<��3�p�RnU���fL�O��B�w5���H�^ {���_���P_�e�.�GB�O��ո�����B�t�P���3-5v��Lm<�A���3E����<s��5(0��-�!Фz��p:9sOf�o<���/5o4EY��_��� ��=�[��G6�Ժ�$��ZgZ�S��w�&3>v@�C77�	�E��]y(��p����G��уBf߯~�����M#�c����uy�E�su4����Q���;�Ҏb�M�^������X.o� PK   ���X�չ�k�  9�  /   images/76cbd0e9-fa13-4be2-a677-68c315f128b4.pngt{XT���� ))" �CH�"��8 ��݂ ҭH(�����C7|�{�{����3��a朽��k�w�����J�~���������@0#��o�ZhA �<c!!�7BBĲ��ƦH,(*A1b�s�.3�7��3r �8	$����s)�g�W_DX}�'*��u�>)}�6�y�H��H�*�[9��V���k�8}g��k�Vz*u�RxX��)A�~<�ƋF �%A;���$!0	b>�$0��=��^���I�;�f�\��"�sエ1U��9��C�D�PA�J�Zv����I$q��I���/9��=��|��Ȑ4�ܲ�C�Ib�N��<HH�Ĕd��l�KB\�]����UQ�=���B�z^�M����@>��;dA��V����Ε�NC�3�*E`�O8��-�"&{�g(������h	�ܬΡNϢ�m-��B��ҭX&���Ȝ!�X�/x���k�ȟON#�^f�8�����F�m�p�+�u�X�jU,���uJ�6����N��ę!���D_\~
�mO�dX�X�r1�[S�m*��1���������L#�3Cb\kw�/Ǆ�֮��O<�B�/0�x�#:��g�S�f|(j�>�E������a%����:	b�-.VYҺ���:w�p����`�8z}�¸r�W�If�I�7xˣBڗX*U�}(!g퉬�E9 /ڀ����#M����cU�
b�4��#�FQYЇ��H/�������yI,�V ��<�b�z�A�B��u����	�S�M�����#�I�ށ����)�s�WXԸSp8/[e�aF���J�}'�B��ۀ�k��&�1�G�L��u��5����8���4EA�+0���}]`�)xCa��"Y�	 ���b��_ТQ��
ᤊ�F}wVD�z`�����w�ۖJ�
u��T4�k�Ƌc�ce[�*���:����a_��:�څдa6�	�/1g3��b�`��I�d ��\x��G����p�#'j��~��4k(ӯ.��z������k����<P9���G�U`L��b.4��]FJ �q|	�����L�t��MF��@��;��W�W��\�띘-�?vAPz��>��ARHHHh���AC�=Hq&,>,)bȱ�"J�I��)J?�E̅w�}PD���rN4�D�R��#2�#���T��@�;��:6��W��V;�:�>WS��'[�G�w�G�c����
e��&�d�-��13�}��ڡУ�f蝺!�����aH/C���";[��0��nj(�$��&�.I_V����8*"��.EqO�F� � ƣ1�e�>VV��RF�
�����E�����쏩�K�G���O���w��WOe���I�T���&k�*sȡ+�|sW�Up�Rh�J+�Y.j���Hq�
����x]J�Ψ�;��[�=�U�%7�ޏ=#7o7�a0o`o(y�yi�s�x�)Gb$}�mso�l�pxx�h�{4{���@�6�����@
Ӌ@�	Ӂ�L���;�{�sX]�
�[���f��2
a� ��#b�3�M��'��L�a�ڕ��@����{�E�Ř�9b$�b��{O�p��W��S��|��J\�6�N����[�Xr\�SlZ�j�o-�-�2�*;-Ѷ�5�ik�Ș��߶��,�=�N�M�ț3���os�w#JGO�Hױi���q�\�v�17�-�HJ��.�&�@���(2�Y�Y�q�p�Wh�k���Y�گV(W���-WZ��1���2kWkT��W�0ƙ���?�V��:�=F<�>r\������ε�.m�%X�ݮ��m\+2�0�?�7q�;��*���rwt�~��At�u��a4C��xj��=x�`���!��(>�2ԾG{�_}s�<���z^�w�+K�à����(u.G�ʩOlm�2Ց �^����;M[�������Szm��]�}�f5��|E����k�J�D�L}&fL�RfN�D�>Gz{���1���n�6˻k�.Z�׭��Z�����^ckb�ci#�z�4&�a��y�:"�3�gy(3��߇&��(�ޑ����_|Z�-�2�ܡ�����/f����Y.�E�0�-�0E1���t4��q��Z�$�FQʺ��u��Z�������vUvf�v���Ds�_�ɬ��t��?�Y|���^O���������-!�����M��UØƩمr]��[9E�c���G"z���3ey����{{{��U�U�_93����͖��U�𥉉�;Iu~�m��\� �=����tw�,��kN�Lm�^��-�m�kþ��S��T����:�J��Ʋj�O]8���YЬД��gr<�+�r��^[[tl�ll�[����of7
W�͉�-�8���ɚSs�H�Iלs���E�QMKʌ��	�ޡ�Jꑍ��r�E�x6:�6�n��������,}�y�~4� ���V��X�(�\n�_�-S2C�֮s��W���*�NV;0q3j����U-�slpěO͚���e��U�T�[Lο�۵�Nwys�Ǔ��8��us�7�Jޛ+���[u{pSs~�y6����ta�L���0L"�������r�j�#��ƾL"4� ���۫��k�#�����Տ�'�jo�'�cRc"�oe��L��g��^��[��<����W�'t�8�3㵼��D���#RP�H��:vpq��� ��|�/s=�9}Gy/ނic(
�8�R��"V0�Ӛ �T4�,�e�����o�U��@;�-�+�׏�I(�����Rϲ9����g8lY�:1߸okU�\��׏���H�.��Ӽ��}�0%Lȵ��7�RR Z����`�7?��cQjЃ��aA� c���A�}���ߟ>���#,������\�<�u3r�K�7o�Ok��杅����G�H�bj6 ���7�yr(pɘ������$�����[}����_��:r�f[=bG3SsnG>ҿ������u��	���,���5���������������!�����ˁ��H���Zr������F`f...0���8�����Vϑ�܆��F~�#�1�6��5�0'��_O��Ζ����9���������m~�p���_�̌L��m�7�-���#�TM��3��으�����J�~��b������+�l �Bf�϶����������@������s���y��}Əl���p�3caE��gXmo꟟�[�ዕ6$z#�R�f'	eFJ�=%�Dq��6\�R!5R����ު<�x6�$&�Wy�Ja|
�N
�T�}�������侫�������9��+�t�}����3�������Hz2�H�@�}	�ar�y�{T�M�O�G��T^�<�u�E#�~|�3QR����\���'48����~(�Ѥ"Zܢ�T�i���q��^8�9��7SP��U�C�KĠ��w7e�%��ں�x�~����-�u3FT�m�'q��υ%�2� ֵ�&��I�������k�1,�5���0g!�߭J2�[ɰ?��#י`!��"+b�y�K�rs�\�Rd��op���(+��s,~s�w;(�(���iX��'l~D-:7�'����P��j�q�'�����c�4��#�ա�C���:?�0ϰizMa??Uj�.��~}�X�=���D�7�҃�7�+W>�T��`�J�0���E�(���H��������L�����I���N�?>e~�֗��n9)����z�r�X7G�U�w�Pj�KMb�w�c$8X��q�sς����TɎ�ģhq��K���hN�x����8\��B\9W��䢑O|̨9q���s<1G�.�_S1d��Ͱn�Ѕ�G��5�h�#���������D��Y�6-j���#��妓E�y�r��1ڴ�E��1Z�q����4CH�;�b*�e��5�0����(6�bLW�Ugy7@l<����T��;���r����V[��i�b��>���ȼ��L2�Sڈ��	PO8W̉Z�r��'`mz ��L'
U�����wi�u�Zё~��\�Jy���֨�ZQڌu7C�j�
��d�/��6C:���t��9�b7�~��ɘdE�0�߂ˢ�J��ޛc���r����@"u�.�����=�lݏ�#�d� �Г�s58�W��?}����`3:����e[�O�?�	\O��n:)��#Df^/L[Գݸ���b|;�9eVB��ڐ��.hԹV�n����I�Kq;��|��Z��4��D���A�Wg��OܯNw%�R�{g�T��d�ܑ�|�lwry�����'@�qh� ��hՖ��O2z��Y%Ġq�������g\�-)(O詇3eb2�.�e#Qꂰ�ā�n�٪%�C	�tp!�ѽ��`����Ov�U��NF}�=�W�Mce5K,F"׭'�0�����)4�?"p�]����AĆ���p�\����~ �`�>x�����cf�-ɺ�����ȴ��Cza�?��%��Z�ъ�s�E����[���7:1�E�b��$� K�!b��B1b8 �!UZ�2V0��d�!P���4~j�����j����9�h�?�� �:�9���7�ظ�Я�ߣV˳Wь��\��iq��U�����Q��p̋Ƴ6����[��q��,��7�o�O��He����Q���]g$�v6��#��B��Hd,[Ep%��g����s��H;����\��D.{]��utR�/4���-&� ���n�ң@�s��DP�iyĉ�9�_)-W�(�&r+� qF�v�`	�%�m8Ɋ�q�ԥ���B$0'������ޘ�,��>�N��5�Vɏv�8t���~�}����>��7๳�?�V:���?s]�s��r3����N��DIb� ەI�&M��f@_��^m�A�G]t��[�3ÍRZ�$��}����l��X�B����L;g���\��W��r�J�I�,з%g�._C�����`���%H������b���b_F��q G�XC�����<�W�����'� ������|	e\�A�߮���+o��닡=�q3\j���Y{�x���[/��7������<�`D !itURA�ޫ|T��A0+���II�ngb�du<KI(9
��xn(uF)n�{�w�&Ze�\���y%���� 貣[�7��uPo��>�xe��6��|�����_펩�����	���d��0�KX$�R���o�N�����ɨ	�D ��j�F��!�a	�M?�l�w��{�О1I�8���׹:5>�슢s�	�ꍼ�g�E�X1�/��ᥔ�wu1s��m
p0��^�:x�'�SL��-���)�\b7�;�8ܫ���K���d�(�ya6�8UbL�q��cv�����5e
�ƿ�v���b\+�y�^ն���y<�	��z��h ٛ�߃��m�2���5 P\K�`w�?�5
�w���u�ҚI��^M#�٠�Ts���0�]�����*�#yZ�v�Gk���+��C���l�J��S�]�K�g�uM3m7��Mt���c�(Z];���0��`C�`q����E�Ӱ�Uʐ�[���� ��-����0�*���!`c"��8햎�2t��� �)n�Z�����0ƞ�9`�L��ޘ}0iD���f�d����$
��붅��<�4�)e�G��F}eڶ�"��H���|.+�������f��1���cA��M���PB�4�tq�L��<-�M� �q��`H_f���p�P��Z*j,޻����
_�U�}N��S;\���A(�p���g��ǃ��x�5���`��k �ᯟsd���?/���}�����1)�Z�.3KP�.�rX��x�(ŌQ���lA�@�VY�{����.����I6�`�C����p������OtXWw7A�߉E[s� �U���y"�|/i���#�λ�~k��N+��d��a���q""��r,�'E!4�J�*V���|�Y\;&l�+|����Ɗ�J��PA�\F����e���k�B� *Xd����.m�7�I��9�چ��_��|(�l��3Ep������*�Ŧ��3�����A���ظ_u������
.��iz��av�9ӄ^9���b@��A-�u+�#Hǩ;F�]i�ε ��/S���5Vu6���TԽ#� �o+
���x�-N�M%�t�!�_���=�n8��j�ܺ�k���;��S��t-�<�.����'�[��yZ���*ZH���*H��q(�_� ����b���e�G<VQ��ot�%߯�����I�00-�.W"S�#��ͨ�=ѧ�qf��
՚��a�l�~C����Z4���}�k��3�-?�2�R3��{ʁ��Y����&�a���v�P�$�3v6�$+~է�ow��u4 
` _2� *� �l�XR�+��/X���y,MOS�o��f�)�d�"���3~WN=!�(ui݆��a�0��:��Ó�(��;M��^�促�I�h`��%�� 1ׯšW�R.���ǚ�9�{6F����K�^L�jb���h�����<���f��^ ���K#~f�!ҌM?�a
��n��[�F�c�H���5��r��}G���  ���F鐅��fW/�S�>�\�i��[%� �Yms��h@���C� V�wNz��72쀚������{�Z�����	��Q��@���ҭA��T��w�����S��U�4��'S��Z<�50敦N��J�8@�?>�{�Md��Յ���KWi)�|{�������Ȟ��	J����Z-�7L�ǰ�Ϩ:�NQ$���O��2GR�<���D_n[�<����[�͒�fa,�{�����M{?�`6��"W���7�C� JX���C^z�UK�S���S)XcA���bU����X�-ǒ��?�*"�)���F��(�.���=��!	pԽԋjጁ�5�E'�&w:Z�S.7����Ŗ l9��hd��p �_��Õ �� 2�9�vB/���(E�"�;@wo��$�B@|qe�J:�2�y�B�Dڷ�8_�~�/y%B͡��P0<����K�O�[/�T��ޏfu��.����s�ZG}���a7���T�?
��Q��c����e6�F@($�1#��l}���e���$$Ed�� ��jZ�ԯ52��{a:�ڒ�&beL��c�9�ݜ�����t b�������	�2
�f��4j1����l����Wo��#t<nF��X+�d��� v�hh�w�Sܟhp�w��	��#��%��yU�ьZ�?.1! ��5�+��Y:p_�C��T�8���u��R��yܹ1�r�5 T�UW��Ȕ0�yKk����ޛS ���}c�fS��E�MY��$c2&`���v�A��5�5���%0��t���y�C�]'P�����?a�Y�<w&�e��PKu�u>Y��?���4���=1RȐ<�08�,��Qvj�o ����m8��:��H�ɋ%��{��u�֌.@/�w�h/�+�؀.p��XR:_Xcs]L>;���ޟ�]��J�V�m�<8�.�	�b`��=�SS�P`��YU,���JG�}7)1��m�U3�=�@�i8=��v�Z�VC�͇R��>�R�X}bZ/F�He������,z��|G���0\�1��<�%8�S'��LǳY�t@�IO����NGf]�z�(HNߏ�1(e)�/�'8��L�Y��tR�p�o���i� $z��K�v��v�v���:'<���N�����HKC_
WNT8�W VD��� �I`��;Aeސ���S|-&r�ϫo �u8%�)d"��l�٪P���hz���V�U� z?�����M���R�'�ee)��i���Q�Q?:/�^� ���v~�X����o��T�7�G�
mt�Q�2lG��1� �)�;F���t(��z���J6����9Pbx���sX�|�~��"�j��:�Tߝ�j�=P_�Dm���+�n��G)T볋V�Ͱ����hͦ�V��>�D�,Aha���B�� ��9 �ܞؗq6����Q�8�жtٯ��޶Q�5 A�������l���B�X�$�N]M��jWT��e�"� cZ���3K��0�M~(<���<�+b�uԍ1QQN�+��#)�ë����x2�gr&�&�3bQ�������J�FܥF���Q�]����@d�A��@G�����eA��y����@$Y����۟m����uH�U��������7�ŧ9/�϶H��M7n.�����p�w�����L�~�x}�Bg��* x� �x������~`M�*E�����〪����Q��*�{�Ր���5�e?d�� ���/;��[�,��^�~�T�u���<�b4�	����Y �m�E�S3G���=���F�����M���'*k��D��u$�2CK,���y��n>�T� ��9g��J��$����?�k��`s��N?��x��a_"M�Lt�������lU���͉|����3�<򌆵����W�B��d�,T�q\��02{fu@���������f.��G r����T�U.}�k�9��9�C��D�T���h�w�.�V��w!�Eݾ@1V#{�C+��\ZQ9'�L)����dI��dk4�j5Z+OC��W'�4_���j��l/��@�S�L��,&���,�z�/g4{��)���˅�N� ��ިW��fVͼMf3�.�[~����tw:�7�k�{h,�� ���w����N�g��.Rd��N�q+�Δ�.D�f�O9
C��9�U�K�����*6�?�Q/zd��u/ٌw��k�듿Ѣ�.�W�|��7��@L�ϗ,Oae�T� ]�C�E� �t�I[�q����t��h�+�ߡ?��X:�w3�>�ڈ`��c�d�_Ǝ�RV�#;qc̓Q�� m� ��/?���l\�K���?�y��L��q9�"�z�1H��=S������S���'�_�C�e��!��	1z��'�������j��C�܋@Ō�bV���s4��8PF� y._�hE�Z����[��SƱ���27G��>ug��������r{[u}�-�]��a7q.ܟ��K��~�dk{��c���U{6Q%�a�adYц��>n�����_F�5L�3�M��]+~�]�:�9[�.�ǵ��4?>�z�i���aUa���q���~�Y��pF�о�� �T��x%���U�;i�|���t�5�sNF�w��qhA�!l0���h�Wu�����|9LH�Ģ�M�E\fTR�|�ڷW��ebɐդϒ������D�	K�&��eu�����1�Z9ry�@[`� ��$8Kpӫ��#S�����2��.��$��ρF����kkr�+.��7��������*T�M^�뒜ӝI��]$͹
Bp�ѯZ�#�΍�ſ-{���*]�h�;{s�#�L��CTK��X=[-��۪��ؐ���q���}�H�D���B.2x:k��ɽ��<*�� ��O#8������fC�8�*\(2Q9�����d�n�<e�c�� v�|�h%�f/&�F��9�7�xw�&����)�>�Fj8y��5�_����w?@��2���Ҕ0o�'=�����,u���ǕN9����\��X�A{�x<�pqe��H#��/6�-�3����W9 ���,^Z�k���MP§���SC<s
��4�4tf�p��_���-����Š����p��<��$���)ve��E�e��~���j�g��`E-����g綿I�0bK]�F_�YZ�����l+	?f{�2g�A�R�n2Q��o���3x��hɟ������Os���`�g׍�ESO堓�߅�	�v_��`�H�w:a0S$�ĭ��i�m�{�Ǒ36Y&�hL�"�u���PpD��V��eLa!뭏*�D�N���2�]�Y�w�����uG�ٷ�IC	�y����p4�bv@F=��>;%���I�ǒ hW�W{���2X���f���9p� z=���\˴Z0# �3��6� g�S�/蓜z���C���f*��ܟ�śU���n�Ƴ��z�������e�+��I"8tD�j�(��l�Ǯ�,!T����������8O#B�yJˎ`V 6Kn,�����Oo��� �2>���1z�ѱY�b��m�UWQ7��k�)��1�2��H���������#������oT�d���&�d�{ȪVU��շ���!��?�R����=)�H����[uE�L��(LQR������ M:�X�e��o����Q�m+�n�d�J8ex�(�Ƙ�E�l�+�}D��"=i��,�<[�0~�����8�U6&
�����׻�@�&�q���Mڂĉ؅I�w?G}z�����<pF�~<P���_5f�4���\�Ɯ��r�Tz�@O���<{�*�T҉�w���� >��w���<��:�Iఐ63
�=���z��Y%ؘI����ab�d�����,W{y�-Hm^��8����Gk�ç^�}Q*".#M�sy�BE5ݹ�c�+W�8������7�����4u���۩�e�'�ضx�A;�G�nOk��@�؜u7�K���Ak�����TrR����T��(˙�����JW4}W�O.pL�ly������1�0�8��7W�f?�;��f����ݰ�~&�:Ű��S��k�#����1~�mɴg���:���*��X$}E�[��Sܧ��4�Z,3�LZ��/׶�Ԯ�)=z���dwo�������� #r�!a7P��e��ea8�����r{�n��@����}�/XY��l�CSn�xq�5Q��C���gH%��ק")�����?7������ދ��<�_vQ��<��FğSk��2X�߭g3&Ve���1�$�����CB��y�H3����DBtfJ7;�9��|WzT����V~��AA7�������w�a�AX��*�V~OY=�����l�hy	��w�Ҭ��KY�ښ�&_$�wR��M*�آ�2{Uی�,�A����5�r���I^�{��zq�ںM�EG����w����m��Qʝ�����~kA�I	Q��y���d��� B� Q�H�����U��X����� ��k��w_�ͯ7�q�3�>��/@&
��ZQ������@Z�uDkt6MON���ռ(?�� -�`@%ғ ��8�Z�k�oi���f�����iЦ�>���_��d^����<��?��B�i"R�	ej�f��� A�c;�}�K�z@��)w|R��5���s��M�I�Y�ʠr����m��&w�=��:�m��>��қ����|`n4sS}{���f��.C/����%�8�����ҽZأE�Ɲ���xY�녵Y����F��wx�XKMzAHM�3u����܌���܄S?�(��λv�[=�3�������N �[:|���=����1R�s12?r��E��t9]
�L6@�%K�eV튡({vZL�f���.�7�����T�\	$��	4>y���ݱ���^{��K����ɸ�x���JĘ�Ė���l�M���jK�<�:�0,�٬\O>RH/B�'�O9l�>���m���u1���	poG�p���H4!����l@a�ؼ���)}�7X�C��{r��_��ʰ��v�r��͂�#����-,@V:#�$Ļ��O�`�iw� ڗ[��%�|�Ji::�Ʊ�6{����2�
�t�@Z�U���df�|>�0�cΑ�BUHr�!�y��>��M$�D��N�2��gsywU%L(�Z)�e~���Y2&�E�iIѐ�f�1a�d,�s��N~��G��?��j��{�U�R-P/^+�IP"�Y|��,�5�I��d� w_�
 m������RүL�<Ƴ�KjK�`n��4��OzO���\8�V�N�F�(-���d -	�&G�X ��������m�����`��jW��r[c�y �
���jL��h��5�Ŝf_8 dM����l��~/@zi�c�?�_�6�U����g�n���B��"֒}�1T��O*'���P~�-Lb�N��Z�$��u�ɀS���@Y�<��+y��$!��1�Q���ܨ�������bΝF���)�Ƥ�l1�C�$/�ȯׇp��xS��Q3��@����k�À.�v%�������]��}Io7�y�-)��%�#�Q�{��UoMi|}�`%9<Ʃ�"ޘ��;�Vipma�?:�^G�N�?PGۥp�d�������?)�V9� ��
����;�"HCJpUv�%`kϝVۚ>�[̉���%7�]���o��+:��!ש��I4�?|v�OƻT�~ں����<��Q�J��W�=��U@��XF�ɪ�8���T;�'��\��`��ޯ4����ݗ�pn�3y?�vI�OݙPX?n;��ny��W[[M��{�չ�+O�km�]�9��$o��t�u��6Ҍe��g�X!	I_��p8���4*�q��D��=ٙ,Ό���<�kumW�^�3��A��~Ͼ�˼�q�,v%���==�z9ƶO쮁�2lt��ۮT�삆C�\L�:v4��,e��O]�hꅳu6�K���:���w{S|�o��I�'���M��x��,	��Xb�^�R�����x����׼3l�q��	�1�y�z���>@f���Sf%�&��C���ݚ@��]k�jĦv�^��j�r�B�"O&�d�x��z���(O�A�="[Cn�e3&�������N�
�iUۗ���}���>�O�z��G� �S��OҤ1 E�ƱpEve��:�_af����F������[�͠Q�2�����-8N����W������V�%����|�&�U��Y� ��%?L$��-�O�smɪ=#\A�OYXf2��Z����oI��d��M�5Zn�X<�~e��_�|�V�A��c>�������O��5�x��pYrJ�{�����k�A;qii�t�#O����A���Z/��W\f���˅�����x��b���)�����*)���p�'� �����,Wه��YaENGki�(�D�8虜I���T�һLZ24f�eQ��F۬�iO����\i��J.L��B(F��q/�:t�.�c�j��,�)�7T���w8�v���qK�>`������>ݝ&�&kn�z�n1_�w�ܛ��d`_����Į�/0�Czz�
�/N�����#Q,d���ہ�a��ּ�g��r�����ǧ���P
�e�G=ۭ.ϯ���Fd���<���U�4����ݚ+�2���-���"��=��x?��Z(����tBv�i��F�@��/��ʜ˾T��L���Xf��5�$�~\�'�/A}�!7���6�<��/��ߏ|_�|M^_���J�Z (ͳ��^i"��B��"��'�SVl}S�p�o�A��6�m�)7���0�z�x��@���:(��J5x�p��(!�w�g����������w�b���I5�-H\Q$�m�/�~�W�~����.�q	i�Bu��������������xXf־U��q��&��U���%�Ieۑ�W�r��$��d�Njq<�ErI����Z~�w�GI k%a%��f��N�:baz�-��#���]��_��q0�Ϫk)3]�|��I>�}��6��i����1�F3 0��o���)ew��w�Iv� 狖`Jm�B���R�'>��"����3m���r�f�`�{�Q�����C��餲�to�ib�)��C���6�ޮ\)Oת+�����%$�Z�\���Jt^��b(�nؽ�ݕkC��hm|s�����!���)��D9m+ͽ����$�c�"	�ԏ%r�|��"�0����?ޅ-j��b�MU���z��9�M���]kZ)�x��z]������]n|���̓qs?�*�u�����pyR�����2�'QkH��G洛io�&\�+)�!t0X3P�D6���4�N �|��qSړ�ѯI`�Z��Ѱ�b����A۪g(Ue�]�ffJ^w���y�k"����L�0�<}�>h�q�?+���6���jCf#��������芷`�������Y~A9�C-]��6�HZ���5eR�Χ��	���˓���Oc
.��V=H8�;��<X�0!�sv�kG���i����xU��Az�vjv_�
ӭ�)���9ٜ��w�W���-Ts&���Kߏg�/���a���0<U� J�EX���W���ۆ)��݊@X�$�Y������s�ηͱs]����O�;a��@��#�����DU��.'�9U��`mv^-;�����ü[y��^�Z����@[�w��倛0�ۉk=�1�]X��yW��8���IO�X���r�K��g��{�uM;�̫:KB����R�n	��![#?2_I0��8��c스�&i�����A/R�<T�19�ߋG\B pZKz�'�d�}��Z��o%��(d�'��d�}1���
�;G24���\ϙ��pR���y��jՉ��1���O��uɨ� �S	6��t��k���K����x~~�r�g,���O,��XKY@)<pиX/]q�ɯt3���!��o������{9�W�@�Q�y[���O0�>	4ɯ�9��&�}�J��j����,A�/�g����'��	�#QA���TP3��J]_5*�( ��6�?w]ل5�ϐIa4J��g�v��	~R��$���1hN����*��.zq�e���	�05�K�T���l�gQaD�Q�qb�/��HŶ5)��`��t]�O�Ҫ�b�S.7�ڕ$���G�-�m��E���x(U��zW�mxz- 7���|&v�%�%�8�*_a wO�ڦ�2���!��l!'[�V� �7R&$��=�*3��U�s@~���a��(���<����tg��*ў}���S�yh��?Wi��KŠ1v��T{���t�x�ʠnݿc�=l;�vx��d�p��_ދw�+/���ƴ�0��A��I����(�X�}�4���F��O�Mc�ӳLN��xAF
��
�0�^�kqSW}��CN�A��]�g���$��c��wl��5I��E����!��e�N�I]�Hؑf�v���(���D��e
dX=k��Z���\G,o����Q �q�'4�����in�	$B�-�JY�4N��KdX���POޣ�B���b�^��)	eտ7hj�� J�~�����C�a�߻(���T�.�L�����S�1!���(���|�*L;�z�}���<-��G7+Ƿ)�;�$�~ʘ���x�?ڲI��VG8������Q=9.�;�������j��aD�t���=��X2���z��^�UE�My~��V��bS�k�$��52���ټG��o�����!���L����mF�����G��yLm	�Lj�}����O�����6;��U��82ml7#s�B�����:�F�u,��� �i��Վ�4�o�*�D����@�b�	�������%#6BHPPsT�Ϗ2�̏\7!����;�F��Q�Ѫww����N���p]�NM��D��z(����^/�踝D�ߥ�Ȋ���D1<!N#�����D��4�ɾ�EB���'kt�w$pby�r>?�*(G�����߰S����譝e�4���=�- �9��$Zba�x-ϧ��*7@�b�J��C�?���c�]��`Ó������~}��+�jw��jW5-`t� X�F�<\��_h6H�RR�b��$n?�,�Yw4CpW $Q�z���Ų��ʂ_]��".ps<<��e-�C61I����ԁ�_��_%W���,�Pa��ɠ^�)C*� �g1{�M@�����-� �t������f���~��~�|9�xJ�m�Pg���ʨ��{�_K�M���j7����oE�~.�����I��g;A�����]
����$tR����k��~�*P���Em���
4w�6�b�a��5�`�.����Ȫͺ7<J�7���«n�=S�ԬG�'���v���8���
���!ÏT"�#z=�C��bv����*�
~�v�Zg����$�L�����ia��|������s7�_7�
$�W���`�փ�s&�a�+Aۺ�"/���|�����F�
����sv�	���ң�D��%j�=��V}��%� �K7G��"ץ-AV�s'"�E��)Ƕ��ߞ�~~�����8��Do��L&��c9��>
Յ��j�96�6\F���Ռ����D4�? O
����y8�����ICX�?�9S7'`�����ΤըJ��&�U���>G��L��͉���)E�ܻ�.��F��W�aU��U�(���7��8��
ɲ_���w;iM�����L>�Of#6D�PMm�bUz��P�)� ���g�fx&�{�U���ĄQb��'}��4��U#����|����Ǎ'� �_��+���>�£>���?M��]4�0����K���.?g�ş���TȪyuw��峔s�z�3[�p�4�.G�〓��F�&c ��F}���.h�8u������K�D��k	�� ���n{L�=B��h�%��'blՍ����~��A|�;
��S&������m��j�!.��no�K�ə���o��M����:� ���ч�����>[,�SX|��Cx�>F��wDfy6��=Qh��߾��,�ɼ��� k���]~����Z�'������~��i
������h��N�	#�
K�*H���>�H2Pn�s�41����h?y��_�l����?�ͯ�|�'�:rTmK�0W��4�91z�5���!�$3b����|��o�kO�WO(�ߴo?|)I!�p�+���C����D?~N�si��LL5X�� ݹd �h��dL ��Ɓ���I��@�P2��4���R2���q�&�y��&�r{XXU���%�������,t.����ή���9��7�xhG+�I�y���x���^��o��r�Ԟ0��c�|X%�UT���d�R����#j�֚�^���E���Q�>�n����t�f��5��,Y>�/����� �fU���V�,�DA 5�P�����'�*��;����02G�I)��ܒO9^nffvk���eX�M�6,������n	��.i6! --�iA%E�S��)%EZ�6R�����;�����|����/q�ff͚��sf͚�ո_�91?���f��~x9����ʪ?��ufǰ䥊�����K�e����0�� �XU���_��E�F����R9�f�0(F6-9��E�LB�,�ë�.O�����6n���'l���p�I5%	Y�dA�]?�ay�Nc�Oo��hOvΘP�����3[�?��۪Xem�B抷� GOp�������%Ŗ�(9��'���06{�A��=��"�̇�|�I�u�Ͼ��V6 ��_��T�-s�--Y���|#x���v3�q����ۚ�����ɑy���K��'��o47�� v���F
u�]�^Ԝ&�"�����"�����N/u���].0�C�nL1y��*h$����T!G>����W�6a���w������4��t;��lA�`�ŗ~.�=m���\�&�?�ȿ�U�B�$�b�ߕ!�0�y{ό�PY~�Ԣǃ�^�R���:�W	���[��4y��W�$�z�8'��z��J�H��Z����=t�0l��J���J
~{�g�)��eV���`�]�}�j���4G�C������{���ND�Zܖ�'3t�eƧ�s���W��z0U8�ܧ�w����?�����@	Hv6�#(l`���p�a=b$`Vs�@�Y{�p���u:=W��~��w0�Mj�o�뀊��~�ŭ>��!�M;��Ñ���8a�Z���[g4�=E�f�P������LG/���Y?3Zc]��'
�� 舳g���z�3�yJ��½�i��3$�}���Z�_�.P]P�������՟�)o���
R�5J'���8����-�/q�T���w6Ϩ�Ϥ���Ӫhy�X,�ų��ܷ���U���8iGB��/a0��O�3h=�L�̨�N��O&~����g����r�u��B�<`��x(4�J�I�F���9�1��x�wՋ������t~F�Gu5�x��>��Y�T�YZ����������
B�d�m����;_c魫q=q�q_B�j���MM��޿��#�1E�9�8c_�<��5:�J"�ʁ0�w�>��� ��+��?}���/������cf�V�N��ڒ�×<F�S��sb�niv���\��9��"홵!�U���D�c��r�[���9'�,�-�C��K-�ny~N��f����}iZ��:����V�s�
�N3^��h��Q�����=�"O�h�����.�̋ˁ�r�T���d-]	w�kf�4+�K��]�9|��п�bn�VD�[Z�UG2�JG�]ͼ�*�00�e�kB��+�n!U���P�Q"����tO�3���h�&y���xk��ը'/��ۤI$v=-{�_J;B�M����o�Z��d�Y}���z؟ȝ�����4��^��}����/�ۙ���H��ȷGW���fg����T��b�4'�6��,=���+�I�tƌ<��T�͡d$Q3Gޖ=�k�	+L�����.���c�L30
�D/��r~����|����s�����_x1�Ϫ0�o,��E�Y�7���c0��� �r]��� �!�t1ml�:s��
w꺗����ɛ��;CP�zJ�(�͏X��ߋ!��Hm�b�������\�?�'��QJ�dz�8�7zx�p�f�I;���䷉w����L~ǔ�<c��X�ɯw �a-��Y�L���}Q�9��#+E�S����c���E���x4$4I���;9�P��r�@��4@�?\���ޘ[��y�MG<���O!)�M��)���+��PBFd\���zb���=-!!t���p���7o��wW�X_�S�3~���J���ۧ4��k$�}�濏���y�`���R���*�bFn�;���$�B�G���E�F�Jr�H��L8x>�����2pyv���fI�ʲ�?�{���fk����x1������?���\��4������w.g�~�Z�,��8���.&X�����;�!Qf�h����(,6��I���Zu��|`��^~)P�i��Bm��	���e:E�	Y��IXy���U;B���B�e	K��j�<�d��{��ƱѲ[�/3���!�	��|å_̶��D>�!�M�����L�"<��R�L��i���W��Y\�A�P���������D`�t� #���J��n�<߳}M	6Ӗp�����=���S��f/g��-����K��ң��8`��w+{�}t��mYZ�C�.�;�R��k�Isvղ_�z�������:��a����_,D|��7��s���������/F���9��	}�3E�����C������
4�N���M[�0NG�/���g�/��1�ӽ ,`$"�|U�	� �����2!�яg&�5!��0��8����W��I�A�eP�w��l�I�4�R�\E<0��[P!�*0P߆�n9�'Jb�#��{��G��L��hdI#�NW�yĳhʄ?ഛ�i��i^΄FS�3�ơNA�雄p���A� :�[w���!9��;�M��!��|�����l��ZU��J_Kunㅂ��l����{x�W��t�BQ��r�4�(_�����Gy�.�C���[?:U�R�������}���Jٟ7ח�[�_'J������z�p�0�����-[������)#I n�yo~|�k=���Ӷ��e�k��O�<�9�&�~xϨ�ߡ?����`���:SR�����A��N+�m1�頱�,���݁J�����d�N�£��ڸ�AN�N���W��9��m�&�;��� @8@�Ũ�a�,Z;a����S$��#	�Rp�8���|�(�����q#�!�M��F&�^������ņW�򀢼Иb�W��:�39B\R��0Oۈ ȀA��m<o8��9dA��/�/h4�0#���@�60Lɮg}�=nnaQ"�(2���Ӕ�s �c���E���F)Υ�Iu���5��ࡏ�[0�b�
Z��A�^b��Ck�p"����gԯXL]�HyBή�����t�m��4����Nh�0���v0�D�{����`ک�W��[9�^q�������D9QS�!��F�5�U�A�ɮ�ނ����F���N�٘@F��ތ��w�����}��1�A����/�ϔ��'(RXw��N��d;5,ݳ�yÊ��%Aύ�M����l���W�hz��$�'�,���C�4�H/?#�~�
r�J��E���uy]bT?�Ew�x@vۚM�Ġ���Uk?�`��(�b�l��@���d�A X�2��TޫxV)��ǋ�ح���rU��*��D	�����Z�z�p<K�x q�E��:(��$��{N���?_��bx���B�7���}����&<��Bc��������f��ɅD�#�� �����\g�|��Tm�t>~�с<g����J�V��)�K��:S{IcԄyy⊁r�ጾgR�J�%��� �&0%}ٞ~���F�'�&E�6�\g��UflB��Qt� �B(+�E�x�$�R9�]^r��Ạ!�a���佤#����Ϲ�j������ŒL�$+w�m�`t^��3 �c/k�1*`C�E7��O6��zP��q�ٙ/����]�lfJ���-3�G��)Rtd�o7�a]��+���[n��ˈ1k����.�(
�,OW�d`"���p��p���bV#|�q��+^�w3h������:���8�=Є�S�0!ߥvB���+����:�����:19�����-���Wz�?)�gt(���7���>����sb�C�`�4�2�"�x4$>����%�Z�V��D.���4k'Pr� PS#�(Y7��g+���$%6=���˕��d��sM��
�4�R'R��1��){3���P�1v��g������f��|Vt�5�Sè��jA��o߉���V2�KE�P�[�b��R��)YE$�9OYp"f˘8��K�3�l
yb�=��K9�j�3
�N˞�X2A���2x��kX� ��wN)��J��o�6���?�_�[��Pѧ[��'<n��f�|� c4�B��M��O=<��qr��bSN�x(rz�r'�qIa��@�^j=ʋ�%A��"��W�}�r���O����]��E
��k�YC>�>��ژ�R�~�}����^�ex��~ _9�GڦO�$R�xą��cy`] ��g6���dG��z�=���q�np(� u��t���o}����I53�ֳ+o��6���������꠴/cx���>�o�tҭ^oSI� ���9k�K�N<ui��,e&�{��%�?�O��;��j���^G�7iF,a�{��=�[~�7��oҶ�pwN��E%ѴS�M��He�V��uf�0;�:s� =��y�1��押n�~�{���������ܓ/~����<���1P��!25��*@D��g����7��2%�c�é�xB�f�׽�f}q������S��A��k:�xz $��q�r��D��*�f��B.�p�Z�����.�1aH���Y��o~6]i��u���	�"�T���4���{�q�FUn;2Ť�^6��C�Ȭ1�!�a�C����T���s�|	�	����4�	�?9�Ȱ<_��(�$�ڱFH�}��)	b�7�F^b]�l:�Wb[�����qC,����k1˄h��H�y~��صXd���Q�#�.[����H�Ä�Mz�>�ۊMb�3��w}8�eT�A���xp�#�Zi����7.R��r�ӧ�k�';�z����#z���:E���m8
;�����Aq��V7r=

t����)mG
c]q0�f�k�f��Edh���ώa���-dk��i$yg�+&���D��͡��9���fs`�G`L���r�a�숙
����%�-AL�o���F�;T`�᳹JDlګ�΂ֈ`�E��Bb��<�84���(��������&�~����/(P��8�GK����m2H����
S+�>�_�x�-2���?S�����v�a�k�9�5��Ə$�9�*1��9����e��$eNKĊ63V��!��0��P�v#�͞��atR�K��Va�"�n	q@یY�����l�� t��&����DN����K*9�mP�/J*�Y�����3�/��x$��Q0��3|��x
���3��p��{�j�?g��Id��~�騁\`�cρS3�o�)p����Cܰ����z�}�K�s]�`!He��a��	�8'F�n0��aC� ��?��w1nD>���ޭ���w�քOoLx��ݯْ_|�~�z�csk�۰5T�K�,��������.7 <����N:�7E��������g�z��B�(��)��U�n�H�/r�&����J�=$7k@���A�~4����#�j�4��k4jP06��ز���P4t�m�)��&�y?�_������֗�F�<�"��U0�(���q�b�|����+鬣���睪�]dv�gk����ы�,D��{"��ŗ(�=&^�"���dJ9q�!'˂|%p�-��T�F�ؾ��#�FoW�[I\øe�޸�6��N[%v[���yl�vϜ�7�LY��j��eH�,����	�/�zWU��c����H�$���t���+6'�1�q�*�����$� ��Xg�>	%�p�|�	�3P����0=K�-5�窚
S��5�����_��];P�f�WcW��ː�{��ޟ���x��s7�^qW��u���<�98��b�ǯ���R�pr�YN��"���~ᯟ��9��#�t���H���'wN�e���>oۗ��$<��x2^%?n�K��N$+�C�����$�M<rS�s� s�f�c���8r��6����=#�`Hn�sڜ��O8�h�}���Z:��u���'��W��vU�����ٽ�eV�i����3g��b��	ǹ&A�oC�oR��5�Y����b��U>��(�p{�'�O/E�<�I�K +����ٖh?:��a:t-��揶5�+N^h�>�v53xjx��5� <ݶ��
0�� ��1�d�����Om������W�����++s�^.�G�T��V�'��f�H��z����l�C��QH�� LC�\Dh�P8����We+��m�p���< pC�B?{���$+э47�eي��j�,bhzX��XY^���"	��zT���:�o�>�(��L��=�&R�؈���NlX윧hsߝ�lL���k"����"�{C��
���eJk�tOy��Ӕ��=�D�gE�>-�º�Ҽ:�Y�mc�"<�o�d�4��r��cq��d�ӜX�n�h��>��JĩR�a��ТwOI��f$���֩��Mw*ˢ��Oj#-���M�Cd�l��	v.�rd�qN�K���o:@���JءG�Wd��'��(�^���/~�A5�;�(��C���4f݄dj7ʎ�b"���^-�J�6i}�{r� ��Ư~��eY���J$�u� .V!���1!KV���ǯS�H=���] ��m`K�ab�w2��p�u���V��z��$s5Jx^�:��2̌:�̽;;l`H�?#���8�N_˳qT�\�7ǎ��nJ���ϠYH��p_��|�w�uh<�wY1tI��\Ym8#
;;#�w�S0�h;:=�-Z��*w�ϐ���z����9�	/*��J���J0r�,5[���ъ�޷�C��.W�0J���M[LT�<��&���5�&m�R�z���D�5>%��p?����I���f��������,���c+�*x0�~���ڜ)ޯo� �<֘;J-�@�B���b�<ۍ&pF^S�A����5+�%Fq�g���ut�޷��ENp߆�@�ޘ���O�,�&�ű�{���5����K��T�C�5�M���!��z�'�k����"��p���m����ݛ��6��d����^��(G�N&@[�ՀyA�+̈́z��ZpF�� _��ǈc�3|2%�	1�W���Q'��@z��ݏ����	�*��._����2W�
2���Zw\u�?'�<�������z4��
7���mE��R#᭱��*��W]�=%Yv{=F����7�����*�hm�����72�[�HV��{\H�h�������y�K�/D��<��9��=?:/��k'�L�&�M�SN��_�9��'�ʶ;�N��hL�=hX��#�Q9��PO�����i�W$�)����87�	)TR����v�*]��.߲��uWK��p6��#,U��i��c�!��̫J&��|Oa���,v�9j g����i�X}�K|� |P��pF/8��E�d/�G �s��:��QØO��썄"�ve?ą��to_U���Qq�S:E{��sF\�y��$����c�[ETNb~� ��?�(1d�3��Ҩ;�%�V��t� #\h�̘���� �I�ár��ܟ�.��S0�5����]�Z��'_��%�M_'I�����-�V�c��>@v��1�A��ܹs{{��	�;��^:j��DX��!�6Z�p
.V��42r���J�6]���#��<
:Xf	Ͽ�A����}��&��������O~��8�����g[�OLN����Mg}A�՞U f@�U�q	�zp���ுHw�uA%�)s�i�˽��'��V�Uu?0B4��@
�~�8�S�s��
'��� �,��Wn������D�	y�n�ߩ��M���l��o����M�H���N�L�;C�l��rfƮ���K~�pP�Nu�zk�1�;��.���})T��&���T�*����Im���rm�u$�\.$� t/
x�5��T0�O/�˳�a���o���$�m��~zZ���VOGL�"�#�N&��}�>�@�����2��PZ��uLSA״��B����̋��2�{��H� �������V�-9��i���M��P����J��<����neoߗPL������v�Hra5�47JS�=�i��Aظ?�Z�Y�������&f��F���S�˔�W��qY��u^�cT�����q�;�p�v���)����2�S�������[���	5�²�+�TDż���V�����h���S�d�5�K�O/~�od��y����q$2�E�jFe�޲� Z��U �>|��	Q%Gd��'o��0�SA��=��9'T>�c�A����=휻��r��i�C?�m�J��nr�c��ţ�O$��G�Ⱥ�w���s��������hڼq�9˖�XM��v�6�A�d'�	m�X��p�h�"�
��+� �u|��,���W�&6i��ϩf�m�x�`��T6�����5�������ˤ�����b��jC���SS*kX��r�:�N���-���:�]�Ou���B�Q��ƶ�B]��˝n>I}O+Ŀ��� �@��&��1�MC�Y��4�����C~�)���|M�w���!���|�d�/Ż����݊�h�ؙk�o�g���,_�<���^���q����.����h�cKw1�@�s��g�ߨ �a�P���6k����J����nz:�%��q�K���A��4�
v.H��OG��0j�o����g�:�����G��)��� ��� })��tF,��/�^?-P�).<_c;�=VJ���w+�T��Q�F�$ڍt/Ӊ����Q�s��E��!����B��c����С���݌�\����D@;�'��1��F�������(�y�{ry�r��ҙ��=g��]_��j˧�{�����o�Q������c�XS�|���I#V��GrM[�#0�6�`tFDb1��T�t������[?!��r�k⹻�~�d�2�p��WO���
oزy��c6z��G� r`��8~��:q]ވ��ぞ�Z�v�/�沢&�i���4�ߗ3�F��3�[j�HM҃�$�����mӮ�,���.��l2���0W|؅�֑F�xM���sd�v_��Du�ME~�AD~��ǃ}|��NPs�b�.=\�=��_��$A��H�B�m��{s����)��������*5���d���	��� ��gq�r��bYȠk>W�蚧f�cc^�.m��!���H[��'P�=�`��Ųq����,�t�#��R�5��X_V���AzH���2�����@!�[J�{��*�t`��JyH&��s���h�Bpa�d�
��&����~��`�7C������Y����xȪ�����N��N'U~�����ʳ��ֳy��4�1���zV�bp�d�a%�M��#\ �s+7��'�F?c�q��*.�O=��	f4W�{�:-�+k=��?�0�41n�go������D1/V�5��p2���[�O�%��:I��<�JC�AX����bH�1�>@R��f�d�5v��2�~=ڽ�}:�B\'�w�Ǫ�����zH��醿Q�M2���\g��xۧ�cԙ�����=�dc����Pi��֞��󏏦��gB�oN�ۊ�������Cǣ�S��zA_.�T�Wnhr��c�yxN��8�r#2�u#�y�����Ƣ]r[A��x���#Ѩ���%�ܚ�Q���en��YEH����mjf�#g���k�(q�IHh���\��q�,���Ձ,�I<��xN��8��Չ-}��ڣ#y�C�����k�_��7D���<��x�mxtﵑZ�b���]���iq?�xi3Dj4����$�M�<y�%�C�E�A�[�}����Lƾ5�ʺG-��^���������<� s&xs��¨ps�g8�D�����e�T������(�ՠ���B*�Px@��eq��	���5_����R)*W˶Fc?s����°H�ز�с�~r��\$���o�f��F=U�8�_��n�h]�bu,z�刖Y7Hz�s N�h+_{
/�%r��bZ9h=3�ֲ�.�=�=[*I{g���_�d��K#������ލH��{�� z�x0k�>Ԃ5U/�k4>i�p.�f/�Dp��0��L_�$c��jI������ixSv=I|g�=�hS��$�$"�Ż�_8�Z�V�`n	��0iQ��V��S���'8��U�����R��	�kP����	�_>�7a���Z	N(��ZpI~���)<�/R������s��$zV��s�iN�&�}焖�{<��/p9�Тi��Sb�S��Y�A%J�L�^�1�x�OПfC����Bo^Xb^�7M��U/V�a�+��� r��tq�c��p�Co��Q���Q�T74�Y!�xf�r������&�|0EP�����}X�L`>�(پ�������x�&G!Ek�� 	7nr$�:�c�g�ΥOh��3�?}JL[�6KR-���p����F�Uע��y�����صV5O1�n��;e��5R|&bS��ݝ����U��T[gg\4�^R��nPYF���~�TE�"&�35xr#.fP��o�$_3������v~�����H=z�gQ �P����� a@D���q��D�$�=4^�m0�"�s�B�TonVB�MY�R��4��_>�6�	 ����u�Kh�/�Qԅ��s�^g���.�2�s�K��Ї�M1܊�v�l����H]Rs��E��:
`�ܹ��	v�W-
�A�PRo>��  ��^滃��wz��.�&`�1� ��輸�v��{[��\(��ς���L���y�O)zg�Z,���f3�����-B�����i����23.B�܋L��L\�	M�a�p��$\˜�{r���]Ժ��Npb5����?U��)-���e��va�l�)6�w�{��݉^����AksG��%�8C����E��/`>`J�'7��F#@Gk{fW����kg:G��a�X�.������d�h�� XTǰ���ƾ� jp� �z����U�Qt�}�)<����:�u�l����j:{���J�S�����:XR0����g?}1:��!3��ڱa#�)&C�@#�):};�O#n� 0�!�4��R���Z@�����Ĕu�W�ӗ��7��O|fXϭ�Q�>k�h���NjZ�	x�d��-�χ�k�	����7o�zL������;`]58~�����9�.������5�	*����J���@8���Ko�0�ա*܅M�,��ь�7-c��V�= a��pF��	z�ѐ8�()C��y�!#�����4�4V#�.����{�sO��t/u�38�c�J}n��,�Oc�.�#꧿`��r׫�ʓ'2|7�Tf�N�E,{"Y�_��\�:�%�f�=�{�%y���Un*�n�o/�gkP���U9��l�r=�"�7]/⇋�\H9u����87�աg�G6��n~���[��/�vsa�5Ui�ԃ��'�\#�������L��������S.+��d�-1� �%4���1�	�锵�0o�蠟w�H�I�/��˯��z��tǽ�s��B���+F�k�(���hm˕C�o0��쌚��g��E���|Ȭ�T1��~�AW�+�)�`�V�[̐_��geź��Oeo�׌�N���<P��i���Ntmu��Y�2�}�/���1��i�B�� �ށ��	.Ǻ�%M�4�i�J$�;Q����4w� ��������wB��e�Iq���4?PО)��Hd�l� `@�<��j��
)�*��֌�����,�]�*>٦;A����$�/�����B��,\�û���0��Hh	������{!��4��9�p�� �5�)c(H��� Oix�&)���9�w�,, j���n!C���͸" ������@�C,���F"q�����[h���H��L��� XR��"��)�&�>m�?:�X��^ ��G���_�=Ql� �/��v�?e;z��'`���@�D"���4�UY�qGB6���[��$v��s�L�P��=p���H���gl�Y��)�i����SKSr1��3@j,���LnLb.���r=]-
b�u����:(DS�J���؍ В]|�����$J�t{�!U��#��m���,W�x�/F��S��R��R7����& �K"�E�{ q�Ș��N�:�b�?����b�����uԹm�_��0�n�\�	8͊���O�qC�+pV���.�����>'��1I:nm�<�9��=��{��Gw�-"8���O�� OˌY�����H4�䯵 g@�IQ�C�V�S�J�� %�:)P�����<�z�3L�nǷ''F�L'R h� �[BY���4��d��V���KaJ��
� �t���W5�a���ʽ	��l��˝���	#g�Oz�jv���wif����+�ϲ�W�k�����GU�󂰻�#r��*�;���/Ԥoˍ+|��g�J�	�O|H��Α[��
�`���$���������×^�0�)�����^5��E� �TM��~�v�{8T��&���%��C�����
�I����Ͽ�@��E (�{����.-��<������\��thF�XE?W�ׂL���w:<Ə��As�2�Y%����+�2t�����R��!���W�C���ާJ\�dȸ����W���[�[D�Td阄�����8=%�_��Kc׀w��H���S��5m�B}�����D�0|��⭥ډ�3����-"���,^������fA���k5ٴHȺ�e�W9.r;u�����i�j�\=����;Z�q� �����!�EM�T]��6p�e�y�/�:�qX0�δ~yrG������i�
��H4Y�C��˃�~`��E5�ֲi�6Z��l�_DCBc	*\����N��v���c9��ȓ�H�:�S������o����T�S=��]�/Gq���/�����Q��v��H��_�nN���.Zaf+��T��*�I� A���`�9u�6���� :��ɞM���cT����u}N�O���OG̀�� �]J�l.TZ�����������v��(�\6�Ƨ�ה�In�?�������0f	��� �e�BTT+vt^� ���W0�rl
L�e93 �%�����ި{��&W�|���k���Vm��f�<��KǊ��T�o��L�N�,c^-5��b*�vf}xgz�̝��w��(rf0L%SR��@J�FfXl�C�|5.�e��������B{�Kb���n6�W�θ�V�RF|�����9�h:A�� �/��Y��"T���B݁Q�u�k���������%ʓG���c�>>�)kVsj�>ŲW�ʯ��k�۟k��������Y�0��7j��	&޼s�OB�O����1s�����H��������ά��$�A�U������*���Wdܯ���ۯ���}>v��^�6cC��A�/�T���Q�X�|9���l�G�Gvc,��-��)G$x�H�s:2�6�l���#�xpC�+�R�c6�d����B"�jJ�I{�4+�d��F�o�,`��f4),e ��E����b�G �/ϤٓϪ�C��m*ջQ5q��K9"�)�������Q�C.�F�@M�dH	�)�8C�`�KK�+�F~�	�1��	ٍ)΍de���m
��?BYS��.��z��P�kO�D܇hJ�>���q	�ҏ62��3���C��r����u�6o�i�G/�����ξM� ��d���{&�(L�P^����`��9��
Ǚ:"��֊�������i���w ��1��$^�]Ҵ+��j���8ٙ��`�?v��d_<���ͨO��ۯָ��eł��w"�5�~eZ}��e�}�]��r�#O�
�o��[M���g7A]<��o�G8ƶ��(�G�Ωf���т�����n^�������K��Í�V�j4�6�X(�5���z���r�;�J��b�O�}�}�jcw�{��<������j�#��ɶUK�e���\���,[������i"��l=M�Xi�C*��OHm�I���W�h#z&������t^�ٗ�oPI�L����nB��{�˿��[��{�=2}(r����La���\&��4l�o�2o�>5r$���ۆ��ƨ�Jո*�Y�R��xB^d;o�w> ׂG�EP����4�~�_f)K4��s<��H�G���޾�Lj�Fk'�M�~0�J����e,�,�Ǐ��x��H�[ �|#�36W9���C�4��N�h��x8���p j�V�B����0�>Q�^�
T}����cڐ���[U�i�%W��9�8���_�����V���N&f�̙��M��x0���!/��H�B��@���C��ƲBR��	_1~���Jέ����G�W;3�ι���������Ng��`r�>x�][M�[1�u�n���Z��{������L�����9�:Ƙ����$������tH�|��Dl�9]%������qJ��(�O�&E"1lg}	����a���~l��p��˝4��!�n��Lt����5�.=c[ϐ�NUq���G�����VY���-9��|��Uv�ˢ��s�M�H�������N�@�%���H���E�xK�&+ǏEPR�����Y�'�?�����q��uV�ӱ��!�O=��Ƞ9�҇>�n\}���,��t�M�|���'lXtPR���t�O���yz��E@�lҭ��W��k��=O�Hg�,���[�ݳ�)8�W$�w������=��q�ҽ��J$�֝����E[Xa 6��-��e��U����V!ڏʒ+�*ʾ��M�cԥ�5-���#YM�J�Q�v-�N�L���c�lt�`P�G���kv�o��E��%�'� �/ʶ0p*~�}�6��&ہ#�Xv��+��?S���n�||"������+�J�� /0ME$� ����W[����+p����5���hH�ȄHdh����4Yj�a߉Tk�l���g+ol��ʪ�dř��kE�!��t���ڀ��@��	�Է��Ҹ�Y��v�r`�ńv+����WL���I����;k�%�X��B�+-Sz"m�l�R�4���~f��^L�z���\M��8��-=��^m�~"�t#^��F���,��
| oB��y�c���بD(?#�t,?ZNK��,���@P=x�v 1U����L�;��8�6�M��o]ᑻ�F�vtez�h�^�.�l;,�,��<U��[b���������������;�ER^��=5���A0;�. ��������y_�Q��c���ђ�}�yǮ�HIV���P;��o~��zpn<�5���d�r�uo�ޫz���b���ӿ���`����Lm!//��
�U��k��$I�zM�y�0�0�����r!�8	����6G�`����0r�Q��1Hf�è�����!�Ο�0f,J1�6�r��_�Tɥ�ms�� �B���'x����~:a�p�
���X+��G��ʲ#����~�tL�{h��'Z��W1�>�9\�����:�)����T~����dm�� �����ɺ��K-]C�����Z�P�Gí3L�{�|�P`�m#��Y��TІ�6z���^�F���^���\@�U�h�~�e�=�pR\ؒԫ����ۨ� ٜ��b]�\|\�懠�wg�'.�z��� ��n��\Y�z{s	h�1���'�!�'Й�����V�M�L�	+�DuN��&�>��TV�̘�PR�1+��^f���T��|On���C��{+%Ց~:��,ݓB�YO�����D�p����w��<���ׯ�-l�����#�۷c����?��}&��Gg�2�N�����؎\�T߀�zw麬���r#���g���:�����Z@�^�h%0�����+�k�Q>���>ӗK(�3u��ſ```�Q̭HZ��g]����.���!P�c�7��@���˕('�㤘
����(5Y����������q��ݛT�m<�ε��}�5T#�h�s*�͹���0o�E}[����sK��e����YA����?��/W�ԅ�H7��۱Ԓ�0�g�J�^����?W_Jd�b*O�s�D��耾j���+SZ��F�p�{�p���.���'��,zh��&��D�mI � _�ק��=� k�l�q�pn��*)���&|rP�;�hEgv?)?:�����rt��B�叢1��='�e�Խ����!eC/�u�Y;������u�zh[~����[&||M�7�3���8s{�y,��G�5�B0hǘ�i�����:��w���:���v�?�t��2y����aQ�Q�����D�����]�e�3�K�夨^.�y�,�hH�GZ���
M��$}, 3�	d���Fb �*Y�J�^� ���0C�h���r�����v�X��$q�j�������ߠ�z��Ga1d}(�@�ӝ̽n���Q�f!س��-_ߧ�³��fKh[͍S�e��yw�?�;Ԉn�W���5�S��F��P)�T�uW���-��`!�b�s���p�f9_<[�8` �zZ�Fc41��$��/}	�����>BN"�\X�8��݋�pKN�*����I���U�ZC7owO�f.��(�N��`ݟn�'I��[��-�D�Gr�&����W\K�D�fϽ/Ŋ�su����l'� ��$3�ڸ���$c���"�6B���������ep -$�������rd����E��~&>-5l4��HY��vF������p����ƎD�q��q]c��(�$e$x�u��7t�(+�%wqTu7���>J�r��4�>$8Ag�u�Q9a��m}��m���#�����>t�Ze&׷�p���U� i�%����Ŭ##�[m��_�z���T�_�vH�c[��#��G�g����s`Ɖ�"�����}�n�qZ#��<Y�c�P�I����p�`nva����^ؖ�LD���3��٬[���)�!�Va�24*t߾��{�s��40H�r�Q(�%?X9U�֥��qJ/�^*�w wn�>�3��/� �;��vT��-�<fL��o�V�;J�e�YC��t���ـ��R�8:�lX�/@��cT�H�`�9�@���(�(�m��2�Q�#�{��hd��B�pG�){���[ꏺB�&�1Q������1��ts�~�]���`^���IrF�@s��������
���ܸ�����*�P4��ҝ������T��p��G1s���tCٮTۦ|�+},㍱��͎�Z���Ak#"�j�����]<&dѨ��� ���|��R�3Lҷ�9��_g����&K$�k���:�K�!(�B�atI�̃h��� o�|���]�#����v�Jf���$�e�deϛ2"�q	׺E�D2���Qf�-{d_%{�B.��yI��;���g���y��x<��y�G9�(�wc%
����S�h-PQF(�ר	�g�n�779Q���L�T��X9�+���b_y4 #���~6>ï�6�9��).Z)e��y��G�ܸ'�B��38��n�bb�+�ȃו!M�� �_Nq-b�Ȱ"��=P�d]�i��45O�=�;�:u��`?5:���P��
��������\�C�d�n��^I����7��ߍLew.�}2lk�#wI~�S�B���IAXh �;8<��d��s���%�)���|_� n��a����N|��C�h��}��I��|"p�]�ļ�3L�P����Z3��Aכ�@T��[g�*��,���%�*��E��Ab3 �'��dH��@����)��gs��iI~t�� �ōAߚ��'����?7�M��}?�l��<g䷔&�b�r��r���=�M`&_�8�fk*��v�ܵ34����8p8	;~���ک(ֱ��̚�5������h�d8'Ǔ
��I�IU�l�ɵ����غ3�4���k^�3`��}]�/��w�	�>q�r5]`����>�w�ݑŊ�UUB݆VL7H-��|���|c���
��[�=Z�)4��GK|��N/%��u�_�z�@o�:�lO;o��i���;�ʂ�>���l�hV��$�ԑC��'�����?���bޓ$,�j"	��Dq5�zQ��ŗ�a3L&��gc�S�
9b�)!,��w_�0e�MAՀ��sA�=��_�q���O[�0��f�mqT]�~�D�ͤ�ϰ�O�Ϯ�p�Qo��_��j!�8I�Y��i��}Y� ��eW�2�����Fr��3lD"C�u���Ff>ҹr󩴻���<��#o�zI�"^�4��s�߇l���7���΍���X6�P��-j��M����M<�� 3v��x'���ﵫ���ۼ��/懦�FU����L� �9��g��8yjO��1��扴��R���L��_������+w<hPr�� �E����+�s�c�q'��Q+6h݉8�.��b�NC�\+�������9�Nڰ�b��J�p��x���� B��Q���P�e�6,���b�E��ɥ�J�a�7~��]���|+��7����ԑ2'����� H��e�v�k�����e���gě،<&�2���9�[x�AA��<@K�#T�j�_5�܅D��C'f2�:W�	!ć�3�d�܉�8#�:8Z���0��wy�w�ؖ�F#d���6���G$K��c/�����2����R������%~M�!ĒL���<�n���NW�t\�9�e.(V`+כ�%E�;.�/R;�u���Vr곗hZ�FS���{�Cp:�	��X���T�aR-�ף�n��#�����Z}��������4J�[����Y��/5/�{溄���f�*�m�.�k��+�G +	��/���p%P.g�ۄ+�*�	���5�,�h�B����f���]Z(�S�T��S�htS�cDI�X|<��H� ����.U�2���t��5��Z�7W|AZ4�p��T-n�>�8p��R����H�-g�I���osA�Ս!!��/�T#jZ�Nn�{�H(վ�]&�UF�ذB.�r�:e��l�v�ۺ~\��؍_F�cY��;^�I\@	$��
R��܄�H_�pת|w��{��#���3�aT��$K��Fo��+��������BR��I0�m��o�;+%�f���O�+nۻe,�*������l>J���K�Z�EQG�t����N�`/ ;.�=���Һ�*�e#�	� ��3����k.�u�1��~�$!��b��@d�o�oZ���	�O�JQ�'f����v�&��'w� [�W��m6�K(gUq���)�#9��_⽣q:��I������R�Ǐ�AȖ�4�C�N�z�r���>ZQ	� �@Q�F���]�T�R�;.o���)J\�����w ;��1�C�WȰ�Q娵n��K3�?��E��LN�f�@$ފt�{��Ѭj�9x�fգ�tDìH���~��Vh��#�������sor����n�c��(���A�m�D�s�$�=IBPR�c�U���V������+C���!��s�%���+����Hd�n��z��#�P�b����B�225n�Df� (
0�M҈��E"��3������ph�ʧ�3�gD��0^~�_3�����L��>�Ī�ɠ��zW�a���y$Mz�N����؉{=h��X6h�٣-�߰����ӛ��
l���F?OƬ5�öЈ�ʘ&?�`3D`Y�I�01��L4����Ra�<��B����l�NK��$a���yȲ���
���I�Go��sTe��3�v}uNJ���@)�SS���!�n���`�Zt2�Y������I����La��>�^��;?W��ʻ	}��M��l
Pi����O�(M�����AD�[N-�C���՘�i�o��5���D�8������X��Oڹ��>�)zO#`����83�8DB�F����l�L���qK�#fGii�xi��70��4}���_M�e�Do�ל���}&|FJq��ߣ'Ek0Q�/2��ء�Jx
k>�t�JW�F�[<J���(��<td[�t��V���~R���7�?���?a��&�\�g����U���L�}>�W/z�i�em�)b�g������$���a-��'E^zȈOz��]��7ž\H�}a[{C�-�>x��ԫ���R��y7��$D)��#~5�,��7�7��[,��b�F��/ �[WL�S�g�FV��*��`�C;����$��G�?�$�>� �������;rT��7���_P�CYy�{sU+ؒh
tgD|_e���n��"B�^��E���D�r����P����|MD$XY���;�����u�V	� 3���N��o���:��W��%���������RQv����7��n��z����?��I�-��hh�rK�c�E��L���7��I��_�\�����TW#�7���	b8"L�ɷ��r=lȭb�đ�SS'!J~{�M�`Bfh@'9?��\t�I�p�V7�0v"x�Ʋ�7��,��D��������vE�5S?F�7G_a�Z�Y~;�:۝�t���U�ž@%pc�vwg`ME��Mƀ��8�j��`�%��_�{����,�j��g���u����Y���T"tgG�G��t���z�k~�������m�8u��16νv��4�<V�:C�H�UE���9�'�w�� �Ba������f�#l_5f��O�Ȉ]8���򽒊��xa�qd �%�n�-؇�Py��J��K#tM�~km�ylJ�+nAw�$D������	�L��w���c"�X!�#�*��N��XUŹ�恇��F�zg�grm�|<af@����C1�7���+�+T &�0$��x3�o:陎to�Q�r
�s������ƞOs�P
�"��گvS�O�l�w��q��AA��E1 ˺P�Z��G�
�ޗ.��J�A�!(ڗo!����-�B]K)Om\����C�mp��A�º_�r!,d����r��Q(���L�i�Qkxߓ�Scظz�����g5G=��1E�~�|>��@����݆n�5�D~��^\(���>��x�%w�JVgD8`�`П��AOo����KG�*��6D2�M��cm|�Ա;[�T�P���ªe�C0���F��W�w��d�7�O��O�lZz_z��D���k��I�@�Sm]�[�}_	'�����Z�Ig � �7Qh������ә�K����W�?���w�����3_붨9̉20^s�[s�n;>6�"D,���?x���φ����V����n �J�K�����zT��"�����
�p�����c�G���j��vk8<I�I��@�jt7a�M���B�'��_b��qҲ�l)d^�ln������7̮�ȝ�,]V�3ߜ�~��|.	�vl��J��䵿�J�f�&o%�rxw)Ǫ�Z����q%��.�=	,���]�yi��DW7���>D�{4|n�캹T/ͭ����J�s-��6�?.-h��Uy�űD3q��p=ڵ��D�O��ݐy1���ǌ;�*�1嶰 y�����`\��1T�pc�f	�S_S�:_�d]x�t�o�'�kV��A��R��%����@.�I�Pd>�_�r/���>�h"�X�+��/�b��2�ph�2�sMϮ�W�H��m�>&_�sY^�R�$n�3by(��9�4`�]�9iC%N
��!��e���r�HaN�Z���A�f�����Rf'�n�C��}t&%���PO��!}==n�P-��Xq�~1�>�8t�Ց�������;�_a������>pg�W�4�Xԩo�����r^:`������a�:��'di�3���VJ{����FR�^CTbH�&�/�y��A�9mo
��+�̀&q��zh���fa��6�]�W�Q3�}����7h��f��g�+�Rlڊ|v�p�����!1^�;۽�<��^���i �`4Z`�kI��L������7z�G�"9y�5�в�y�3�B�ņ�:�����xD���/ϰ\��Ǣ��M9�|��o��e���;[Z��%�
X��Z1u'+F?_]:Qq�(���we|���D*i�V�0��CR��[iY""�T��ތ$�g�S�5�$��Xo���,O&K�=e�}�����
暼4���y����{w����EtP��M�{M�ay�A?��5?��{��~��P�H�3�$�X�g�0S7���%��V;��5�j	E�\,�}�`^xIx�DW����n��x4���#�GeK5n��~�3B���s���I����i�#�����/�dl�!�[�f*�_��,L�oU1p-5o�	�Px���P��"��]��ґ����y,~����>%�����ʘ7��բr���F����RѼ���yh��upUx������OS4���ؘY���1���M8;�sd���¹�>�@�k�Ԋ�n�.ށt���%l_���e_hK8ɋl(֧�$�h�5�֓0�=u�#w�A��bKaCi'��x@�{jy�'����pi�l��{W@��t����CDpu���7v�:.�S��|;��9ߧ�63�L:Ǣ$�m��YN�Exc�`��*��dM�f-ε�E [���gY��?��/}��`���Y����B����>�2��$��a��w�9��8"��� �5��=��^�����k�h�I�#"[(��ᡣI��!����W�W6g3b/�t ���%�����+�p������H�R� ���&�!
�C�Z�t�%��R�1�1�Lrym�3�������l��@��b�M�esƲ�ǭ����b�������F�1b�
e���e�=�����E�P��(^�=YZ��w�g�W�7_va����S��{�ۤ�sK,�Ξ��^xg���G@��[Sȱ?�*J�~����`���M�����P�����+�>C���2d@�vӏ�A��W�y�0�V��wҢ�o��K���C�_���T���=��ӯ�B�x�ҥ�!w�p�0v�{�:P�D�-D=��^�;���~g�l�hj����S���<>N�|�����9�ؾj�����|
_��-EϗXC��D��{���FVw��f]6�=��>J.�7� ˹�<V�˧�kx#c  ��ִ�W͇By�ҪFY�G���e�R��e�����&���#�X�V~��s�,F��|�I�i�&=�2�����>�0�P�֚�����J!�ڢ�E�DB��-J&o�7�EV��ѡ,sY( <W�nՉ����O%��Z���ҩ������/w����-�I#v�Rd)��	��`�=�^�=_"�(�K���)~��m$@�M��X��X���n�����Z��5�׊/2��+�2�RGX�.V�Q��~R޹�F����h&���_�i�n�v�ߠ��j�w��N�`/86���  �Rb������!O 5ޥW.N�sF�K��ߘNv�&V�jY��k1�dg����������f��Mm|����bp�,1��2I��T^�c�H��+?�_&
��RB�V�`Ys���$��$���� ;�Fo_Zɧ>U��]+<�Ō�`y�=�d�{� z��c�w�8g����#m�����CyV1�d��v�<=����X��c�'����X%�W��gޫ�?R"���iy-d�v���-�O7�����?������S?�þ)~��Q���V����ű�MY)}�<G�E��~*(o�r�y$ό���	B)��J"p˻������Q^�T��5�3�F!3X^d_�M_z��I/G�b:��^<T%�=Pz̻���	�J�gݞ"+a7a�4\[UX��v�j��#?���w6���u�n��|���B����Ih�zz`Pߵ��~�v�j<8N+�ҘO�1�9&�H���,�𿦲��f2l����3����S�.S�r;"\�L�� &7v
���4����K����A�����٫��j:b��������4������9���������i�^��Ժ�3i�����c��m�%Gd�Q�V�Z��/�D���Qu<��L�t}��_����M�(�F�x��z.�c?�oQ����ɷh���O4�h�%��-��i�Ix�W-�S/�dQ��}��4-�]���M/C+�ֿ5q2Q�}q7����+���&D��g�8A���@J�9�9��B��6�=`��U�.5FꜧX{44�V5.R�11����,]�*I�QQ�s����2�w�Z�~$�g�YyC*+��2�yDt@_��r��O�T���Թ4r���Pv�^@R��q8���WvP7�̱O��/��B-��_�sJ���0�
��HkcyL}��Vci�[�w�E�+���NCMN_Vz���q~�$��S�����x͝^�0��\�	|�ζ�k��8	F�3�$���[�(����B�m�*�g��Ƅ~�<�� fImd��6��@��HNR8Y��@F�{^�S1�Q;U�X� 9v%�|�	=���ō��Qc���_�7=
����Ã:��xst���#��%��Yh
�����#f���6��}�FM�ehO5��`,��y�E1�fq��u�z�R��5�l����^��J��B��ĩVʚ������ח��̷���ʕ�H���~��!���`�����X"�� �$ǽeLp+�(5d�nq@�䰽<����6��u�����ޑ��T���@㜢�l��S�_�������A��e M�����X�a`����L����M�ok�0��U<f��Fz�z�r-�Ӟ��=��+��W�Bp�u��{~�Gۓ��ҟ����5�/->�Q�Ӿ���$����)��+@���t���������Od�ӧd󪿢嗡�L��;.�FD���)�'���^�R���r�~~�ͳ��R�ϒ�z���;No���j@�θ���=)�����l
�[K�}"WX�����O�/\��hy�C�L�1zM�}�n�����^圄c��9F?��_�,� ܶ ~+xi���3�2	�Υf��1���G�E�*���Z���;�R���Ǭ\�JЗ��ݜ��~�Q����A�wT8�����h��	���=���e��0�����k��GM�u�e��9����\'l|�L�F��ޯ�I���<��x��7�({�Z9 �y��\:�����e~|��2n�e�qza�����9�2������n*5�2بv�Qd��B���؞$��Ax�������I5���Ξ���_�tj�PHl��[���1$�e�J+X?�p�p�1��^ƬBM�ϰ���WS$&��G"삧���MZ	f�^S�=�'�͌��*L~�����Ԋ 5���uˢƿL����Xԉ��wԃ<v�jxqƥrt�������u�{Dk=�l���IxE�����;�(|��ئ7�fcP�Aa^�ӏ��2)7����`�����k�.gD�l3�D�	��� B5&��ĈA�s`�w�|�؞����*�К��#����&9�<߇T��	5����U�7�B�q�E�?�v-\\�+��~��)��V�S+T���?PK   ���Xd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   ���Xb��O  �W  /   images/92294c6c-e025-4a92-b2dc-6de1496811f5.png�u\T_�?�!�""�H�J+ �t-!�t� ��t,-R�"�Kw�t�����Q�����=�=>�{��{Μ93sf޳w�׊/�q(qPPP�e^I*��������c��쉋�����KH�����m31��������9N�s��!��'�/�>	E��l)��{(����%��m�s>�C��~��@5f��@F&��An���h�oNN��iϕz�ED��r������c��\��'1��R��Gv�R�R�6�(�`�{P(8�J.�4v�(9wg]�\?��$GyB4��+ȇ1?�1�V�7��u���ʓ2b0\��/��Z��>�����o����k��*��C'��|��$Z>\����8�^NV�)��#���$�R[v���Ŭa�����r�HW�������͵�r�� ��z�p�\�u%������j\�+�D�=�#kAn�W�"ؾr�@�}��L[��T{��1V�������p�ѢG,���J3��_0.�58�F��X�+�j����v)�,"�gz=��r�&�>��������m�Q#���˞?3����9��}JI�d*�6xulBOn����yl灶��殄�3���>"i#�X.ƻ�Y;O��>����|�����%��}1��h����KK��\˃^t��jyѢ�eU��^"9���*�;E����z�*��ˉ���ਾ܇!�/����/Ð���s�*z�N|�&��(�|ǌz/1ι��$Ӈ��^n�i���.���.q�{B}b_zjɀ'aO30�$��H%��	�	qҾ>xBK���	�:�������b��r}�9T5��/���V��}e��#>�s-`�6O��B���f�����嬺׀>��}��I8�	E�,4 -�����)�t�i����7U�ow�y|���>����QN�m}8�L�^}�D�9P�PNl�m��Mm4h���z��U��7g'�qA!/���|��b]���ǋ��Q�o����Տ
��b�1[j����-h6��wQ*	���9c���m��/�M>1�#J	5����̥,0c�{�2>���h|���7,�Z~>z����� ����>e�r3ڻ���',n�'��������Jy���}�Ȳ�G�i��#�#g�;��P	�'>��.|��X�wTf{|W	Եd����7�0��uq.�u.�G�'E�2�&���{�Vڋ"A�b���b��o��b�~�f���<�{�f_WS�U���.ۏ�i��p�����Y����<ᚒ"�[i!,,Oǟ��BY�Y��)_K�P=)����dMQ�~{U'n�j����q�������S�E���ڛ�|Y���
�ӹg�&id�[_5k'����q�qqɓ�O�i�����{iԫxjK�4�Id+-���*@��%���ɟ�,�ɡ�V0�I^��e���U��ϛUP�U��_ط=�<�9�=�1h��/7��Ѻ�=b5H388p0�5�7��U�/{�yugx�/~�<f�g6�1l�Ep�s{K����r{Vc̓E�LAn�BK��J���Wؒ���%7 `#���=d*�e����ǳ&�ǭ���5��W�����5B�4i�B��TːňR�b�aK���S���2]ش�ek�P ̾/k6�pV;^�}��T�4V8c=��+����I�$K��Գ��_%��̿�����ټ����h�(�X��(����Na7b�̯�OXէm���@a3�T�V#�8�PMc��6y�©[�U4�[�����+`#�
z۾���u����w��dE`�Qޚ7L���Q?XZд\b1f$z$j�Yx�!���rw��R�����Z�*4fD�a����飃z�� �7�ϻw�1Ep+�z�R?������ֈ �o���ٵ9<\]N$�Y����l'�޼{㛳l����_݃�v�Q�Z�����4�BX�T����/�V�M|�m��YΩǏ�(���&��� �c�˳�~ak��~�i�Ŋm�m�-�^�^�������b�}��$w~I|�/�*�22+�1�Jy��������G�Ѫ�C�C��9����V򛬢�E�`=_��d�z��dd*>XX��.!)� I<�U���|Qv�>�6�]]��h{N�u�c_͘�Ն��J��\y����@������籡���ƇޫBE;�8Ƹ�0<�x��h/����G���N��Y���QUFBY�7�бy?�4x�5UQ��4I��c�h{uz���F#�?��,���u�lڿvvR���I�#��W}D��L���s����q&[j~�T}�A���93�.����������4�o��1�����!v��vK��~IY�~#�참�f�����:+�O�z��Ɯ���j�R�5�)��/����AT�W�u'�+3�̓��J�)#b��xK��C�i����g}��S�#+�ZA*]qzo7�s�S�̃IhQ^���{;t��|��Z�֊�R���iUV�v^���rr��78m�,����[OL[n�m	�m��l�P��g�5l��f���:sLC���B=wLz��g��\5,y޹��
?�8�n� ��43"����%��^t�T�־?��o��~�DG`�{�|u;a�h��[�<��%�ꐺ��p<h>6-6�����ѵE�h���y�=���ɗ��ɂ�YO�A����EG`a�}��bj�i��'�{����*P�ޗ�
���#���w���ٛH����hS��B��C�|�P~��ǹI�F�F����3�m��cOmE���D�0�>�ܿulB���"_�}�Ŧ�ĕ��kC��B�d�q貗T�e9��5�kj�	I�M �~�jȘ((�<�X(訔(@8DQ����Q��ܹm������������_؟����D�`-b�p����7���;ۨ�7Þ�H�� g#;(����@�(���m�
b��B�ts��(?�����j8h(���8�a�P+����]����������^�E�ᶇ о�b����`! ��^f��� s�Dq����M�%����0�98��@�����0;S��� ���bz�ۻZ;��[�3�G�/I�������9̚�滁!��A���O������b�?3Y��Y�@��'��������]��Is+@f��ܜ\ ����H������������j'�n;�������7�
����b���(�0��Dq*��R5R�K*�g�?f�O����Qk��Mp���|�ꂺ9��H�tٶ7�P!<�WY��+�{}Pў��?r@����W]N�4��\�2::	�^�;����u��)���٫k�����m�{��q���q�i��H�c����2��(��D�7���}!Y)w}Pа�o>�0�I®�N;3��G[���S�jf�İ�l���Rӥ��V�B,��<�[j�X�=zt\�J��@��y�䋑i֟f7���!r<����'��,��_���[��z��c��g������hI��:��a.��u�$v�n}�P����p�Rg����a+g��d���v�N��N=���¨T��5�߯:�qϔ
"�q��U+�\����D ���� g%�+=X�
�5��k��qXc��uv�����sg"\iɒ�c�6A�U��{X�Lチ�[�33P�'vloN���l8�.7�q��ИӃ��Hz3����%>Z�]�K�#�K#F c�������\�4:��P{uy���c�[���~Lb"[��q���֡�?b�}��:Y�^�6x2N���W`p���}}^ⴥ� ����6}�R�NU�V�ȁ�V��bAmX|Ӓ�w7x��V�[��gd��o����C@߄�r�	�9�Ѭ�Nbճ�)��~;8�NZ�*�/w�~΄�~�#E��>
o$C�?.9@�{����YQ�Y��Q_���)�g�@�]��fF�c%y�~��5-�>Xȫ�<f<�mJ�w�7F�K�]�:���}>�����*�t��&��������@s:]~���@�p��H�x����ST�դl�v5�k~���@4�F���3�b;Ӥ���k�ԻW�����CK�D��R��v�3lo�Vos��]F1N�GV�$}��g��.t=�{����K]��;����?qL�d^���ץr4�6�a�t{}����F���G�Ǌ���GuqO )��6�v��k?P#�����
/���g9u'���K�;lB�o��#����«=L��4y�e��~}y��`G�4�\-���Ȕ�se@�b��S=�k�N�����xzޗ�K:�V��<O�M{�0�=��Siq֞_'��״]ϥzu����1MzY����6A��.�!r4ѫ#�C+��&y	�	C�$����dm���!�$#�Q��p�g��%8&�x�yw�9���D� Oh����.Ew�+�IҢ��zn�G`"ح�3S�^�Ӎa�j%z3��g%��}�<���� o�i���W�%Qbw��囙'&���}��L��\��ܳ�m��z�C�ɾ:�#IBΚ�'�9�#�nH����K�z�
�i��>Cտ;$׌�b��8��T!�7��b���bgW�z��5dډ�bc<�d���KIQ�r�]��uL�W'+a�W��kfU��c �~��Y�ƾ�Ǽ�Ic��_�}t}����Ms����]拁{w�����O�\xc��R���מ����l�+ē�)��oO�.]����d�����K�y9�s�٪2.��B�ڌ�8^��~q=P�+�F*w��-E|��՝{���X�oqS�����H�Z�hq{[ʻ�y�]j�MS�{W�m{��'ԇ ��[��R_q�n<���{W��u��#%��* E��q�uaB�!2�FI�ς�x�oE�ǯ�7�x_��@J2f�����o�������~% =|����ʝ�]b����[:���Ru�f���y��Ԩ��_��>��Ξ�L%�V�G���{�8O57���yb�1�u�m/3�S��9b C�%\O��|�r���Z��|����� Rn2��!.멪����d�������d�9����g�<���Bu�Vd����\cկ���"���F��P�e�ԉ����]w�F�p�߫w?�k���`����7�Üژ�} �׍���۩?�m����E����S�����a{J�ˡ�������xN���y�Q�=�tq�xm�H�G 2��`����[���_W�v�oe��|HE%K>�v����-A�j��f�5�lzSf��#Cn6����|��F�a�>��}�[,�!lL"�������j��QY
	�eddX�����y�`3��E!������B0����h# +�4����g���e:���Ϭ���6��s���w,8�*�~��Ri����Г�x!�B"��d����� �H����s7A�{��<��.5�"U�� ,�X)9Q��ȿ�����˿l{��r�F����^�R ittF��t7 �E�ܐ��v��V�#Q�~���׬�*)6��q�Ͻ�4�����- ����?�||��Z�(�ه�m�Z���峂d!8���]�qV��_��I����&U~��S���<VS���rU���?�U��O�x�)���8�\:�_�QO���q������+�ج0eʦ/��eD��
�ROҤ�F9i]yÍ��Þ�����)/V��ȁ����y�W����ڙ�O�Ҫe�Mm1K�����݃���F�ŤwQ�����g\6�2=��0�GiBē���~ˤ� ��5}�"�BC�43�W2���K����Q�E���*{�7�`iܧ�C�x�QL ��դ������]�P��x3%;>�_[x������͔_b�1m�d�;�%0帴\�?�y �x@��Q����������`��fq�?����3�����Nn��>�x��\��*���ÍѮ&9��x�߿�H�5U�y,oMV��ŧ<)�@F�sg�<<�ϖɈ5<��iE4���_�YKW_�D&�Z��S���� �A��+v�T�+�v2]��I��`\�_u�qX;���,���4�󌚚��{�뺘��Zqm�:j�|s�v�0ޑ�<��6"��,��5�yƕ�A�l�0�Ɨn�8�(m��z)� �}�ⷑm���
��Z��X0FoZ|�IC�(g~�+n�8v\
�B��m%��/Ъ��d+8R���$����a����U��6���ES�^��[Z�<Q��\���蘴�|A�LP��gR�N z�}�!-^���[�-:����{���w����]m��~� ��	$����Oګ�R��y�R��:6����}�[�/��E
kn�Mbq(♸e�4d�f[O��:Üm��D�@���6=�?;��k�]
�3�My4�'̎�8k���{�ĈwL��Jq���!˟g��S�59��{��[�7 <s$�shJ �.��AI���� �s��6�$G$M0ޟ�aӽ�Hh��5��\���~$�r�kW�c.���2�,�*��"�26zʌ�/ &�£��:����S�ZtɛG�(�S�����,߂3���+xSs)C��H;.��#�ƭ����G& ��k�L����s�ֻ{�.s�U���i�K&T�LԞl�D�B�P�x��Nƺ�q�B)zu�2)`���Z���Ӝ�F��{_��LV�nL���A��5���������W�q}Q����K<���5{���6q��E�R����%# T�Tjҽ/hW�_m�|����e_�(l��T�X+1|���O��Iud�E�&U�/&�*�io��O��~&8)�bEA^�0Ƶ�[�[�z��[%җ����W�G�I(�n�ʏ�?""��sE�jپ ������!����@�uO ���G]�s� �,��q7u��xTŗ���a������g�J���!G��� �e�ޣ�ç���M��YI��"��NY*�=7��yo����-��'�x�<��k��7O�u�&�)�q�� ��ޝX>����d�Ec���Ufby�M�뻀f��'J���5@v%��x�4
��3�lE���,!+[����Ӹ����q�t�y#2WL�]��/{��
�]��Cy���o]]�ӥ���9P��{�u����Ƌ�������1���[�F�/��n(���%LG�6X?�����gd��J5��g~�A2�%�aʮ�1�����R8�]V�"i#���뛞Fvc<�h�
�'�	��q�{�&�t'E-��\�=�Oԋt<H��K� �7�� �N�����~w�#��L[�{��g��~
APA���ɃX�^L�!n�KX|~�sS���?�a�>��i��.V�s*���Y�Q[��[V��` W�c�#��W�S�	�G)���8l�q=��nC)�p�2�?�t�X���sU6!����!q��*\�b�!����̡�7��E�H��L"F sV.|����7��ے�<;��Lz-��	�J�.��K-m
1�ךFr�H �.��U8C��S�+c�6��/G�oB�H�V}g"�O9�����&O��A�ge0����=���)�_2����V����G��d�;D�/���g��@8}c��c=�P_wy4)ڦ��H��1hW�A�Bb9t�$�ty˸#�I��A�	!c��p�c���'�.�.�w�_�9.h�ϬxB�83B-䔿��sW���!��ɯnye6�?E����$�0��|0%�����&*�,��U`Z�[�&t�ʖ1�D<��|!n���ARMj�|�[Ħt�{ }u��أ~��d����}�T��W���)'x�	^Z��ȕ΁�X�]��[��'��2��$O�[dM!��"�/��ҝ�2���E�$�ŭ'C�H������,��⹒���;��l#cM�;�m����y�4�נ�����]��#� "�l8�'D�.D���N������8zA�Jr�"�ߐ/7l'�eڝ�h>d�p��ϕ�ʇ�>�cW�������J�k��?(���So��w�\���&P�ӻm����_�z.��Ţ[Wu�3K'���_.OZ��a3�'@*	��>�˻�%�o��
N�%�2����I)ܢ0!�K���`"�!�W�Ȥ�.��?���2��@��?��r�����ꛮ��N���� @<�4�����/,;�� a�K��	Y�@��dJA2O�.�{�����g��;s�7nH`z���N�=z����ˡ�K�k�u�]h2��4��i��/��ç�=�ݏ�G<��I�ȿ��*/MZ�o�-"O��7��ùϡ���vKEM|F*ݦZ�au|3��#�p]A����GI�­f��8��r/��p�b����N,��J�~Ԋ.͓L�L\��p�gLg���Y5�}:�_Y�S���7�CApZp��3�mD���W�F�E���yŬ��;���E�����n��[�]����nE�y�vg?mY~I��B,��(HѨ����P���I�y����Emd9��pf��ʼj_.]�n�e��vT����x�Y��[�]'=������~e�^�����+�I@i3}�{S۫�$��]=�,;sz*>�{�FM�M ��܍K̇���$d=z/t7�F�y���⍚����6�� �Y�4yӥ:- _�Կrr��Q�9�	������S��|������p�5l�`�z��m���6����~���p�O-�\�MNx�J\�K�2�/���c���)Sr9�^�{ڪ6�d��,N�f/��,M�
Ky�-�����*?��#fv� �4�qj<����(>p@��r]�g/^�Ϊ�Ԧ����8#���12`t��+8Y��{z�2�H̃��q�F��j�	w�mK]<<>w��^�<ͫ��u��*�ݓߜ��A	w���H�d��h�e��=_�c��An^���Ml��T�R@k�����������hr���츷��22��f�����F��܊v�@}��N�A�5�QVS���o�>��W�q�v���~qo#�5�QcKX�)?�����O���Ew�H��y��/���Ys�2\z��"H�F13ҋ����5n[%�$������쥃�kP�ٴ~�r�쎗�F��d��km�.�8"����	��
$yl���Λ;tY�RȦ���QNMR�8���Z���ci�1� ������\�Q��;����.@����w��'Tp����J���mR�ț��r���?nT���X;):,�= #�JH�ll���8�����C�
�ٿ�;/�k��n�ӧ�a��\&"TD��U�=��Sn���g��#�ji�����)E���++u��ғa��ѯ����}M��bAP��҄���� ����r��N�`���;߼ӱ#�ϿH�MC���6ȼ;&��7�N�Xn܁��d0t��S��Q"���l��o��*�p$��y�����S8��u�E��/V=���<�s��ް���AS뫿<�"і��t��4$$���r�P���8 }4 7�QM0>�ٴ���ק��3�r���O\��� T)<��j62�8�(���w���g:/y��x<�yAIM�B����}����6�Rs��l{Њ��L�y�C���5赿���v�ch��"�u9�7�Z8�-����P���=;�aX&� ��-C���v4L���E�b`��	����Y)��G�_To%&L[�2������o|V������n.��V��*�����9۵�������Qr!01�Hk�ݠ��`��s�Pe�_U�:���~���H��r�`p�;�r�މz��R�kI�D ̤W4����b'�U�Qv*�>�6��^LpLc�*�.�H�WL�2���TW��2a�@��;��vS7��B$qv����ޢ�3�aW�%_��61k�;a��O׻���+�8�϶���zu{��w������h��t�  �^�G� �Y�q��P�?�of5L8E�'\��m�s��ś��ߜ�r^��'i��B��g�Tb�O��u���ޜ9�5_3t���G�MC����?�,�hՄѹ빲z�H;էV�z���P,��Z>�cx+�=�Ye�3J�'K�4�6���&xX�ĺأ�����ٺ�H��]d���
 ��j�rq�C�^��.(���K�e��:,n�[�ƅWY�Y�!��1�8����~�H���D�n��:�xnh�dY^��<{5�.�����󓛨�^�&���ysޠb�aV҈��y��7��Xe���Z��`1���ݪ��%�y�'W�j�z5.�>;�Z"�ݲle^Q�Ƣ�R6��#����:��R�s�t�^�D��`j�W�П���gJ^�b���9��Rٸݶ����L�����֬+����q��&2�tW�9�!6_gv? ��\ƚ���R�Y?_/�Y��S�<�RQ/��Q�N����3��8�w��nr�u�ps��e�|QT��A���B)a���L:�)���:�R�FuPm�)=2����Tof�<�fM�^�>lK���~�d'C�ȭ�=b�u��,���(ѶQ�z�$DL�,x�ϧ�u�'�&N���LϪ
ϴ�:,��ꝩD�y���0Sݚ�RuOV1�oHv���f��ed���A.�:J�(~&k�J����NL�0e��1�,�J��k��$N"��̳��H�
�������~����eXE8����{�NU�wU͕��g�\��F{kY���ְ_��E��S�7>KT�ҪŤ)@�e��6Z'�nbK#X�RW{Yhl�;�=S1|�*�zJrU�)���T�i��Xn��U�q��G �4��q�>_�4xc�,M�*<p�u��Vt�0��y�!��zx���Uk-��*Җ�����a���YnwO�W�R
7�bj��t��u
o"1�BG`��#!ح�Vi�F�,i~� X�jw �~�i�6}P�R��1ãt�4�*�ኪ�?��P�������bb�z�}������\��� M6!f�`�'{����?F��^͇{D���)}'wۅ�.��+�;�?qZ,����M�W*r�	E#�M��^��O�����=�-ZשzF�-#�i���0�_hP/�Y����}��~�`����LQ�X�N������g�A��x�d�c�'F�Gؽ���M����Cׁk��Z�gGI�İ��7�/3H�A0����Y"T�w[�7��&萬���&��@ݜ���8x ��f��"�-g�+hғ���^�!���P�����G|N��|�e����N�������@�  �3UA5�~-����\�>/�ڄ���{�8yfl�&�Y����><ɋ��;t�$�uZ~��_��5��y�p�[6���
ld�g=��=��8|`�yɉ?&����؎�KE ���Ժ	&�)����������_�u���"�@nA�����1��"�.p�KY�p.�� �ᚸ��QG�$�|kb[�_^
p�5Y��=��~�ew�C��JN��i�-��oܶ���S�R��H�Ƹ ͒\*�L�%f?'����E���pr,�%���O�����Mu��46�d)�m����!�k�0R_m4_t_~���Uh�}��>��b�}�7�CU%
��6B�s/���ܓ�����$��帴'��j+C�m�ǯ'K�m�*�׿=l�y���-���9�
�+�:�-/���=�R�H&�g,U�W&M#X:i�*z�4��g���e\�}:>Z�t���7���#s����	qy���ht���[Z��e������3@t���Uٛ�^��8Vs��r;��I��\�Nr�x���Oy׆�w�VvN���x�ڦ��R�{l%��^�O\ݙR�F�v-%:m�fC)Y��X���ˑ�z'+�i�G��u7^�緡�4�ʹ�N+{�r�fl�l�6G}��� �Լ���R_��Y��E�[�|�1Y��sN�/(N�Q���up��%[��k!4Z�>�j�+dcs��(���渾��&63��e���Mg�c�z�dy=��P���;�4L�ޞ��\���f6I�8�KIW���	���!�f2��u��T�;��}9�O���y�;�#�N��ݼ������f�>���v�޿,��dW�Q��6��D�q��A�ǬD��룿\��Iy>%,�u��lE�lI-nQ�Q��3�q�� �E��Avor���"l��=C���B�����fP�����
9(X��(x��(����
�L# �x�]z�B��'7��?�(�uB��vZ%F�֮�_0�0JI�L�����V�Mf�a�	[�3,d�<}V��hA���Y.�U�B�y���5������
�A!7+�0Y����������y����N�S�ӹ (����}�ή��¦� J�L���4jŋ�»��9��M��򑚤飠Y.��:r�r��)���6.�sD��r��������R��龩gM��:���<V|���Wj2��|���~����ϣ�-8�cV��p�d�+�Z<q7i����z*��/Bf��u��L^��v`��7.�W�
�}�������Eə7��6|
�']�i�l�k��:W�7���M,�٢r-h�6��4=[�+�M陏�T?��|2���ߘ��7v�\�q,�oT��*�CW�a/$N	�Ί�ֻ���WIÒ`�����1rz�xei���DOxWQy}�052iJ|_Q���d�
-�U=\He��|!�'>1���V�
�*`>UJ&�|N){�%�-A1Q2�b��\�M�I���#won�����󶉞�wq������N0�T��!S.�l�PoV?�P�ct�<�IǬ� ��[�_�"B�F�׼.N���o�R��<�?�7s]H�eW�Z�'��hR�:�zwƛ����9��}w��Ʋ~���B�K���w���t^u]���B�$�5%(H ����7��"Ƌ=�p���G����B���qF1��a�\RˍbU���p�G�'r`���
���ߥ�����6���W�^�B]v�  �6h��"3�m�&�ꙇ��WR'�� ��m�e�Q��KWl�Ѹvɱ�����iM���A;N&�9���43L�K�����;�|��b�Dc� p�3��c-4�ʁ��%��x���Q�>��!!�V;a��A�&������q3�H��oS2�)VDr���7���$b��^+�-�YÓ�&&�ދT��aŭ���P �\˕����[掫 ȓ$��K�:o��͟�j`HLL�I���E�F�+�������X_��%^/lj�&�A9�O�mMhr��(�@.�&�z�!2R�i�5Nz0e�|��_�ص��]:b��t-k�S�� =p��o�1��b�;�}����u���m��mg|c��T�M�V�8�;����ٌ��7���1Ic�y流�俵�'!􂐝� ��{Y������� .��|I��I&�M������PS/�ܨ�n^��1��[�CV��v6x����ƷG6�!ЈY.���D	YSl�`��qN�Z����-'s��/v�03�t��j�t�2 ic����љ4G�Ո�k�\��Z43��N�,��|��l��,�6�U�5W�=��Rw�$vjU.��4�=�p��\*���L#���eHe�>'��Y(H{I3�ܭ��TfAx2�\;s\�_v��݉���=����{k�x��6�3xg�h�H�h�H���#�f�X�.�ˏQ�į�ݒZC�;>���A2�5Ӛ���Ϯu�¹n��������|W����� 9/�&��ֲ9lT_�gE��Ia��=�̄hP����YU��3W�p�����E��	�wԱs=�l��2��bĐ�j�lW���B����J�����-��h
��>��hf�g�Q���Vz���Ox���R�����B}!8a�?qo'1���'[��u��D��H�l�X�ߘ)߅ނ�68"�bQq���r���&%F׸�܆77��k�,�<ӛ�'t��)���U�z��L�74�ے<�YF�:�)��{:sBM��j����{o����	�TZ�!�������u�0�V!����@wQ{�5X�4<�{�̪>��1R��V&��Ƣ�y]g[|T����v�v���T�z�A�L~\f�V��Y����}�R�롛�LT��Z�l�׹��M=�Cޝ��x,�b�����G��o�����@��RU<���-�v�Ꮞ���V^,J�O�������ُ�����]O,P<�h�4x׌ Y���"\ވ:����VF��]ZI��<$��V�&�~j9�^�u�m2�u<�� i��b���L��ͭ8}���x_ȻD�C@O�R��ؒk'O �~�ǝ��t#�J��G��r��-i��Hv�~�"n=	���$��3��j�B�"�M�N����b��!��G:�bU�Y~E���Q�IY�ū�������"Ӯ�3�\nk(�n�T��L�2���}Q��0P��O�L�{�DF<S�C���1�W�^ڗ\R�Uj��癠���Q�0�K�����>�iВ�"܂���^q�{�V��q
�S�)2�}��H}*�׊\d��6���[���	>����C�p��D�I/�L��K_����G(����%��3���avɑ�}��_�-�9\D�����"�x�4"bfb�wR�����{��IlI�>&l��8F��=�¼�\P�kو��y6���U��]�-H��C�Q^�K� �#�$8�#21�t�J9o�DFژ;0p�_�F�m���:Ӊ9���~�2��[�:0>�H�rg���������)h�Un�G��ȵ]~��fc�\�g�|w�����s����wV3n|(�>��o��e�!�͝��1�d���J������Y"�_��G�ǹ�c���ź�ǚ� ��^s�6G���e�<��pj/��@k�_H��N�.�Ǯ���U&�Fƶ[_Y%a��]Lr7zw�mUo\st�&Y׈:`4��2J ��`�$���%<�b)걳aRGɪb�؃vf�/��aCg���\�����G��,=�lT����:}�1f6�eE7(X�]��jo�;��w�3�g�Ir�S��݁��cK�/�ks�a�yz:���ҕ�ȷ�1�:4Z�ݭY��}����*��_n��6Jߩ1��땥�ͼ"�����Kd�vҋ�Ȼ&�PW\T�e���f ��9�,\�[�?FC���3nJS��$�r�;�k���&׏��8�3�>2]ҡN�6w�qg/.�޿
�Ke�	
-ﲦ�s����]�V��8��R��ac���e!��Wk�>5�w|�1��LC���V�o��&�D
Q��	4>t���V�����* g�^����9 ��D����K�Bn���3`� QϫU���7D�C�� M�>�@�-�� ��+��X{D�Ѓ�77�g������m w!o���W�wS�'�$�y���r�j7�	q�E�Cl��s[9D�g�o%Xc��t��) �!�nx�Of �EH˵ܲ0�;��k�^�7+� Kdv�s ��d�������Hn$��K}SS5g0U�KX/܅=�p[[�T̝i 5LIZx���>�6	=����//
X�������o �<!���tm��BySQ,Jg�o�\���_i"�q d�U� N��/�72�y���O�L�\���Y��:�q�(�4w�?b�,"��8t��ݎ�V���1a�|�{��̰4��x����V_�\hY�lV��)�������J��M�$�/?z����V@N+z���r�%�CG���o��-Fc(y�ed1�X�6m�lST����m�I���~c��,O}��$�F��?"EL/��p~�:ތC��ݪr�q��s��u5�r���ڙ>��4wɻj>����x��e���������=��au�������Τ`F�������GG��$m:�G���|j�0��B�0����L����)��Z������Iv�b�R���VL2�y���37�����f.}�HU�����Q���a~�3LC��5��aZN;3"��]��ņRq��5�P(S��{˝3�����a
�jdXD_n_�z���y��b�����;��iRAFm!��i���e�C��z��uEuuu�Q�MMv����嫉 rk+7����;׽-LC�R�ۍ��FXI�|Xd9��3�ၻ]î?2�&��6�����39Ⱥ*)����3C&��p}8`�,�b��4��s�dܷ7ƛ�3�=�G�!�6
k{v�2�v���Ϸk���j.�]���a���j�iu1��8�
�YA�=��WF�Շ
���Ff*ffъ��$ӡz�Ϯ>����a�11����n1��iBgr�!����c8��i�a�G��=�	,)��d�,p�J���h�L�5:��խ�'V��r+ap�HH�m=ro��(�l鹵b��K%5����c�}n�qV5�<�X��NR�X�ѧd�NHs ~������H�]u5k�9��v��y�.��Y���@E�[nVWbi���u������g\Wh������W��=��JBڡ��۟؜��P�qM���9'kN�ؐ�J���3𡄗���e�B�;O���Aq\PY*7\��oo���f��	7=�WU�/t�g���ݥ���~��B�([\��*�0�G�ل��E.�4�z(��1Wa8�0~�*^���Q���/ݴ�,���{;��U�b����3g��d��y�jJ�#�����©לX�@�罹���`�N+=I��n�a�^#M�ؕ'.F�.�?^b�d	�{�MPq<	�����镜��T���B*b13�:�?�(铅]���8;��>P@%�)CA#��e�V-a<#kLH��k!��}}n��qS��9V���Uj��S+�h¤�ce]�/�1A��ܭ֕:����-���`�%d\ݏ��ۏ��u�6��.E5�7k��8�2��f�}�G��C��j_�����?��ͫ}�Ɉ��ε�3��������TBarW�E������&���1�D���s�6ҖsN��a�9f�Cw,�BV9��_m����������}?�������z}��1�e�����K���ա��5Y`�mĲp�d{�T�<(4~g�kѥ��L4��t"�{2�u��׬��1|e��E�D�ԯ�nG�R�
�G!ͼ�����k6��0�5ӄ���v)v�=X]6�#�����7�$͘7���q��5�&��E�AGY"^�$G5a�Ű��+�).!�Go�z�6��k�8&��.{����u��IĚ��;Z���w��-����>���tuuu?���!�$�4��o�{�=�Ŝ�{a�"i��s��Gp~�*����^�q���[�+�3�u�Uti�惗(�Zv�-Kܩ��wT���I9�?s��]$�Ɲ�v����n���Mv-換�|�YQpʹ'F���c�3�	=o `�E#ˌ�5V��W�lr�
�!�t�9��1[&�g��I`-�X�P�f:���l�r5{�O�8t���eǩ���\W4 �W_�N��������1�[��%���R��LӇ�z؄�?/o^C���Vqcyp�(|�R/����8�̵d�BgY�v�bT�C��K?CBB�$(�ϵ�vi�[�p�����K�媉�c��kU.��gv��w?:6��d�l-�f��+���fL�k{��'�<�zv"9)�{��EN0ğ_�P�a�}����^��F`˝m]u�+��J��b���G/��F&;��ǎ���	/k_=��±/}��)/��Lt�i��q���~W�T���[����Z�+�
�/@�=��8�[�Cr�b|$�X?T���x*��`g�oC���-�o-����KAg;����i�nJ�\�O�!I@�aN�yVT|�MC8�kd���"�����2����;bݵ~��BD�m?fG�-��*�C�0�ĕF�-��ؘ�IALI�.��L����1����1�_�m�6΀?A��}:��b� zh}[ �Md�g�|�'.dW��35a�!��P�gXf��J�S�&4��]�μ�_�o�V�h:�J����_��Ʊ�Y�a��A A�2�ɞ�]�G���T��%��ø�,XIP��CVf"�ۼ��u������GǪ>f���xv�.=�����Y��i���^�ԃ+�M�4�I�@�?�n��:	�[`���x~��n�bz����܏3呋��`�c+�\��F��#65�,����,^�E��Fb� �1.�p#@�~e9�T�^�)�8� �[Wm�S $è��슠RQ��i�����V�7\(�4�F���*-k<�Wp\�O������3l:ب&���&�F!"�pB--����`�Yr|#x�]�Ѽ�4kMD���I�h-��m���*M���������S�}q��S�si@������uTA��b��S}�]�T�*�e���@�7�%����+��Cä�rzU9fPESA�A�\+,�T�h@G�O���a���3P ��*����Oƃ�w��<�`gkb�|%��ή�~��KS���d����%j�N�:����mi�JUy�	w'5�� ��T�l��ԇ�C&7��DP�\ۄ���SֿdJ�Ա�6���x	���i�:D�.]���[>����Y��&Є�3q�v	e�"��R>�-۷��+���ş�yQ$��q�!)	߆�<��67��_������C
��&r��{20��|��[����)���F���S�[nB�YH
���S�(B'���M�ԑ.�2��#��ܨіa�����.>u�(�(�w�u����0�k��jH���
���	a*�n~O�Dy䦹ڪ��	�	�|Ak5=b��H�b���ˑ��F}�|U@�Q�V�Ή��NAN[�#�a�b׹�4�P�%w���iZ�I��7;�*/�|�~)[�0�^ǥ\]��怨�uX�n�����;���y����n�Պ��b�
B����O1u��,���qc���B���D���Ed��{d�.������@:d���N��0sb_,r2����n�
���kV#F!Z����8F)57q$P���k��5��c��N�
myn�*t�ݚ�Tt 7Md���N�Fh���7��ۍ�}��q�ͧ��󇤠kQ�3��]�O���?�g���8t#�6>��%{���ۢO	,��
6X�Ćm��(`w�0w�j<���s{/rq��އ�S��=��^�6���-��聼�$SB�ȳ�:�V�ٱ �w5j@]��O�^I�М��C�P>���d䯵�"��DV����Z���9�g��CY�:��޼�3�͖��͏�W�&��#.^��i~��	���ȿ��.,>k�N�4N�qSD�&�W���?r�F���y���$���s�x��ض���|���A�<�dIm�zw22tA�K=�t�UbiI���ک�C�p$�@P[�t��M`;\��s�q�YhsJ�)���E+d����"������#y�� �Z|�o��*n�{Sی��)ݴ�pX`����`��j�\�R������K�[���q�d��r]��=�;�����m7}o��l�V�TT�j
�S���z�?�Ge����.�!��a��(+j2�6�_A���/=/a�7ǹ�8��3ſ����N�dM�����Jv����P��ǎ+��?��
�~���Ox!)G���Y^������C�Ԑ����Pr$X\����Vo>�<s��$��D��� ��n������u�ZƬA~"�1����Q����=�m���̄O��%(��Y�w9&�t���|���u�:DaN��-r��e~�ց ��c��C	��t�gS�O����]*���ur���g��_��t���x������;��eN��Ђk'�ga�6t��Xx��
C��#;����97�sİ�����[E�Fdvת�u�]hwύ�r�3ּZ�ޣ#W�|���p�XO�r' Ȝ��ϝ��1 {}g�E�i�,��>���^�r=w����S�r�{�d���x㸃*(���&�#-��,�|��fr��AUͽV�d@V��:���^���ן�u����-�=�;�l���+٧�r1$�/J���廉e�+��U��|4��p����b��_�M~�  ��"{�m��۬�ꘕ���3q�PK   ���X�^>1�5  6:  /   images/9756906e-dfd1-435b-853c-fa5dc8217a1c.pngͻwT�M�/�&�
*HS�N�Б"��"(�)$��K�ETz�P$4��H��Q��J�p�����}��u׺�J�=3��6�睶�
--�S}�H"��@d�4T���X���C7����!Sչ�x3P����h�
�9pE|X�(�^����7�5A��q1������9����2�������A��׿=�*������0�����{�R=@e������T���A腕�K������>���K��/{G7i/�;[Hפ��;��#d�hhs(9��8ą������rpp<p��K�<z�ow�N������4���)�	rr�ߗ����ED��nގ�/��8�!�t��,]m��m�9H�/^:y��޹�o����e��#9���,`�`��}!a���M"Oz*�m��7|d� �Cr_���}���4�����E�kO��s��n0W%'ൻ�J������0����?l��g9���-39�Z��H�Y���g^���34=��6�F��趠�����`��<�?j���cRb��I��#� ϳ��9t\|�C]��)�V�t��������r�r7�-����f��I���j��%B���� ��3=`�K�ρ@�oci༼�U�[�Q�G��H����$gg��Bv`W�e�lO*$>9�� ��c��۷����>(�[u�3��^�{����I�X�f����A
�|M�B�q��$�
N��e��6�!ק����d���n��+�.</�K����v'�k���4 \��)0�Ý��G�m�ɣ�k�%��X�	�nQ���u����z7k۱�"IU�TMe�l9S�W��`hA
x2�(v=Q��Ý����Dޫ+1�����43xt���7@ �8�U��C�/'�(�Qk��	��vK��`�p�������פ��Ȭߨ8=9�.|����ʕBL�� n�pj9�%��(��(__�����xQcT�uB�X�$-h�;5�$W^:�C�'���ã�������r߰�>h��C�JL�����Ϣ� ������)���F>�xlJ,S����~��8X���sd���!����f'=�w�����X��yv�	�41����؊G�?V�Q���q8u�nΪZ�6 iq>�w��m�;�t�ѱ�r��[���i����x�����ִgv�;�t�*Og�9���i�̨Α�O�t��]���K������ۄ��%�����:���^T;o'�M����	iw�[�%�{KC���ȝ�Ic��2��!��^�_Ӛ��r�r���
��0��Vp��+��-X��轕��7X������/�����Ύv4���̇F9�Z\���]��g��=�T�=�Z;�� �w�SW_]Ԅ�+���ٶa�rͻOq�eu��ZC0K(��Qk���Tm��V�[0�]�T�]�x	0�yu|1�O���Y����r�G�D�=7,�5��1&�$�o�>�F�Q�ձ�m�FZ8- 7��L=3�J\�`Ƞ��
�̐H��Ք��Ϙ���'�%\b~�n�.��I�:]f����j8x�X\kXO��.}c5��>?��a����zJ���a멾&� ��z����������7Y��f]���>IK�~�F�-���A�.:���a��9����V6�����.K��+,h���Br�����D	�%*�)���n�/��NQ1xuϖވ�e��?��]#W���]폳���(�5���狹��5`ߢ��<�,����=$�a�_~s����F%P	�v)�������U�D����)i������r^<Q]��/w���龥�d㤘uZ�{Y��cH*�.p>���Ul��y6b5����
/�)��$U��8� ��+�iv�Ҳ�V��I�2��z�}S�ΪXb�Ҏ��M�z�I,?��H
jT���bϔ�\Vg����N��l��
�2�6z�<�L�Bh⒨���Qv���T���.�B�}s+��(�v]}L�D��v!��޴�Ws���)o!���������Sѻ -����AF(��ZԲ~��'C�;�|"��}�{��b���UD���KQf>��o����r�ؼ��q���@n�Q���b��W��f�m�2� �	f�~�F�*Ѣ��=�G�-+]�{ֱ�Hz�� ��j�p8�F=Lr�E���h�mB�ea�E�w�� 
j,���x���h���r�&^K0S����&p�	�� ��8�L+�v��~�����ڧ�KcB b2Q�X��û��T4n�wo�ڏ�:T���/�M6��9�{� ���{�����y�y�IM�҇3�I,`P�*\���O�t��/ �����<X�΀��լA�|-����1_��� ��2ӆ��s�uN`��0!G�ڸu��V�����xm�ɷ��M����bm�ة�#^18����=4����%��O91{�Ůwpa�E�ǲ��e���9��,�E"����ɤ@���hv{ټ��C
������BR�{�ȌX�-����Z�x,���Y�3_���~'0�U�)'ٵS&9�� �|��݋��-ۣG}� M� ���B���!e���w�8z��?�P�w5��}D$k����o�<H�#�+���-�^Y @��
p�#S��0�Ϸ�+ڠ	�3H�J�K���.���*���'�W���de��Z�<�6��hA���S�)X%^b�T.y��0�`��:��O&�Q���5�\0�n1���˺��>d��|E(r8��|�ж�G0�sO�̔V5��Y1%Z�:�^TM{�yVi
��o	BZ5����>��I�x��
�&�~M���?�����Ç�@$�=3C	�9;a�j����3N��XT�T�im���no��XX����jIEs���|'._�KJjt��� �ڗ%���x¬����,�{4���|6�R���S�l�#{𴽅��@r�����}�J�x�->R�,|
f�䷧Ƽ}KSq��g��哒1r\��M�����6~/6����]�|���^��aѳ�xɇjj�7�+2
������6 � o����ջ ��b�����T\V�� t��m�����S=�0���J;o��+�8�27RV7�W�Wo���&;G5+	#�;�Z�P��|O��C���a�v��3iLD��t��r��%�A9S�3����Xwb<E��)ry�wU,��z<��ѓձ���r���Gk����.x�E� B�x�A8Z�P��M�jp����q/�uʋO�a��P"ɗPѱXA5���o���nWB3��\���+�h	q� 
��n�5�d��d@�$,t��h&	��� '�cVk�d�*�C\�Z�|@�������2�*7� ��&�3�HΔC ����U�_m�K�К/=դ�Nd<��a���0;�$��y� **��8��e+�*N�^�׫0˜� `pT/�Q0��> �����䯀�Wҷ^=��K4=f�Ɖ���b�e�������ټ���q��]�<�{�YzN�� б���=?���=������ �In�bm�"��D�?���� ���Y��yJ	��wJ.ى2�5z�GH���r�ee��W��m�߂�u%������*`���D�6�]I��eg~���O�b��AH7퐙>�8V��aX5ͨW��'N_��s�{�Ώ��6v$"#����g}��g�Z��sN�i�%���jﾡ�p���ÑDs���&%�?goX�Y�)g�=.$@�&�G]XfG�����/LI��@����d�̣*�ۘ+=�-����/�Y�Ug�I��m���'P�(����XM��\��梜Ąs�3 �7�%&κ�&�`3���+9��Z�@����A����=���N��=)�?��;����6���0�]�ߘj�����/r���6TL�k]���%��a�q���@|�� ό9k!�;||]s#@�D~j��N�O֞s�	~�ϰɻ�����"��^ �*�u�/;d�{7(VF(�bv�����A�����������r:��i���՗�LV�ib�rꅛR)����)@W��L��怠�j���Ϊu��~ޕ>�7Ue�Ƞ򃗺��]I���,�����³S}��&̩�{s�O�]گ��]ŊO΁,��ch뾚��B���u�P TRu\��mܛ�5���S��4y"3�=��eHa�5;��h�(������I=��1&K��,Y_5�ۤ T��h�Gk�&���1lR: ]��0���' ��G;�rRx���}�J�)�=�Y�2�=oΠrc�o>��d��+)p�IC�.N55|��v���O77�dɎ/�A�y��p��Q K>/A
�?$����$��\��U�m��c��I��d6����3S�ރ�:?"F�wQQI�����b50�H��*:�lZ��XϵJ�6��>C��I[c����sz��[U�(.���kq᧩�v���6OG�[XHL�WF	��v�[D�����BYE�Ҹ�uT��H%��]"+��qK@�����|�_�Z^ �K聠dNL� ��=��P� �xdފ���]�
Rܿ��'�i���0���{A�ܟkk�7����c��6о>��g&�x�.Ơ��k�w��S�����ѷ��"���?}�|ӷ���D�T��}���k�o�������<�>2��1�B{)^���kOup`���`W�
s��f^���
ጣH��3u2��P�/��B�yK�_��O����_<��e
�n��:ލ7k��,Ԫ�LTKMw��<�.��$��J�T�T�X��;G��k��Vk(s��};�9S��=t�&
/�1���������S���t5�Ck)��\U�9ǫec�5#�Mާ�x����b��=i&���ℤ0˗����dL`�s�@)y�V��n�g�|�f,�D���I=��������wf�Z���ټ��[$��hV����􃣍@{�i6v����"�5S^<�n��-c���cRzr��p�ա ��R��L90�j��Cv��z�y�^����'���.:�?��2g�ָ��s&~s�|T�6#�]��ַ���6<���hƷ�I�x&�ٽ��eg�G��^_��Q@�vr�al�fw�ٙ��|����K]����R]sG��\{o��YjPN�żu����lê��wg��]�Ӻ"j ��p�?������w��΀Bc;�v�}�Fh
ȉtY�|
K5�V�QN�È�8u��7�0Yl�y���4��tI/l�-ϝ��[I�#�5�/v{p�Nqa�L)�
���KJ�4��V3!�����j=��n
���<X����	Dhf[$�9g�@�⡌�S���!�F�J˵E>@�f�D��-y'W��S��6�L�;��]��8T'�Y̫�dys�d�9��ߘ��zSU��au>;�_~�~��y������{T������� ߬q۞H�ʅ�w�l���n�>F<؂X~�F�3$����O �͐� �����bPT�oӵ
C����Ms���&w��Qߓ�� �s�=Z|�u')�����6LK���Z��ӫ1�>S;�"�C�Q�y��wOBHQ�����c{���O)��Ǥ��h�x4Y[1�ata���3��qb����_�;2��KG/��iJTY9�<��ɍa?�;�?��#�,#ٌ�	�I	������_HC\�Ŏ�+=���:8�[��j�`�k;/Y�?t�z�n�_ho�����{��=n�i��|���T��~z�@hɼhT��WO��F*��oc�N���y�o���������+�n�l�.�9��k�1�KW ��й-}rA9�fva���H��s�0��Lz�˺f�ڝ���ʏ���oD��$���Z�lg�,��ۻ�ǉǧK[�c���|�N?h@���f?¡��<K�a�\A��o<q�E�o*&4,���X�S(�<�I�IxY����:vr����5��j����`v�d�9�Y�_�- �o��t"wI���s��'l�}=.E�$���q�@ٓ�1}M�����
�ۃy1S�/(T_6���'U��ceZe����'��J�_#mO����e��V��Z( ���@�U�\ө��G�6��D�>89p+���h@��xJ���䟣�]�%�Q��Ǖ�ي��N0��2���ъ�<���� ��E�� �yX0��q�xD��)H?�y{"��׋�T�G���^���r�ǃ���y��u��+J8�|��Ih�"03H֭�,�e�G�>{b�2.=)�$t�;,�<U
�ഺ����oW6P�ZJG����,p�|�gs���\�7��.�}4���%��eUDdK+��WlOq������VP����� �huZ[��a��L��F�?"����V2�F7�����wyS��f�U���]�g?bN�C���팤҈�ǝ-�A���ԦF�m*'���}E��g�ճ,����HU��S�l~��;���#ޣ4Nm��9�/���bW3o7=q9�l�"�Л���:�p�;m/dO3���ZV/ӾN�ZP�;��t��mA�q���2��l,^n����l��n�~���j�٩�_���MG�,�I:}Jo���g-�I�%���%j>P���;��t��nzz�I�=���K�t�l���:Z>}f�L}�Q�Z�[$���{�Y���r�=���c�U�Rj���h���f�x�%�\e|�t�g*ܯ,�g
�k�<��?�a��>�tM�P�5ـ�[`�a�j��P!��ް�Q���U5'�rkg�kNř��A��7�AW�h��z�2��Z	5МM��8��k��̖�q7s˟#CՔ����_�}�2�Wb1����e�*�
3��i�s�����ԩW�Ԙ�})cy౗ǽ-�}���&8Sn_(ف1�>X��bo���~SpiKgs)���3� 3���ܯ��ow2\Իp�Q��S_�$z��O���Vh�҃Kp�cs��D%�<-�l0sύ�0��y?x�f����2��Z�8�O�gƢ�m;y�ֻ�<�Su�}�IQ�f���3G<��S��þu����NX��ogi�������ȸ���o+���G��F�ܔG5�aY]��r�CRE�DS)1�7l��ԧ�mÍo�>��1m��,A�{�}���x�Tt�Pu��MU�0���z\�3��B��d���]�^�=�I��F���7@�=��:8�g��5�I�qB%�P��L m�Sk������S\�^~�ru���Sa���,����O��b�m����v�L��w������;�Npu�s�tH��#lz� gя���ߎ%��W��]��f,^'7��/��Kr��2�{��sp0�>�]��ZW{�̄��G�V��&{J�Wl����9�:�t��@r�ฤ*��q\Ca��Nm|}��/�6Y���y~�W�j�6C�c�CS�#5:��P*���dz+�b�̽ݎE�@5�d3�B�yF��{0�T���ޏ�;;���ў���o;�� x<�(��:�zr�Ob�u�]h~A:#����`�4���g��;���
�2��U"�����HX��Κ�b,<���� +d`�?M<}�Ͷ�&%���>�iN0
b?��v�#����`D4��ԍ��T�Z������lܥ��(�°(])7%��{+�z�y�f�[����t�bgd�};��)4ߙo�'�8=�a��@���"N��B�&N�vj�����ûr�,�"����?~��te��>[}y��=�����m���S�	��׾	��KD@A�4�O��_���������v�^[9�X��l�zwҹm2G2�{,��DT���e�|�2#��e��o�
Nt��l"#�t�'�
�Wzf�h����@����'�t��ؘ�R�z�n���jǖE[�)���φ&ES5-��M?�%�.7���%�Rr�O�V��������e�',7=zM�F�<���R�2�-��#�g��}ᑡ���UC���O��m��,$��2 ����^�3�J�c�f)E�ײ?�i�?����|b-o��a�Qt)�����OE��x���1�)Cl'��+Zt5�~����OaF�t�m0�nk���<B��ex�N�ר+������g3)	�I�	]w�2U�I�n����X�[Ъ�{;[1��E(���������5�Gg'n%Q����Ć�y�����k�ݧ_>��]s�yo�{����{/C��J�%�2�ERN�cmqϳue�|zn3t�-�z%�\|�����ﺰ�Y��2�֋��u�m"�3��?Ȯr�Ut���AE��͒���nA���+"#˛5J��uƻ��2܆�㏹�`��
��.G6��R��I;�^��V,��b�H���z�$�{�OZſ���ޟ�BۧG�E]"^3�	G/��[�j�{�S�]τ��/8���*BQ?6���`��Ɖň���̙���|���+���
����"ӉL({*�qYVj ��A�����%8���B�[n�ƋS���)JH�+��!��-��T��5���g�x����A�� *H�@s����m|֎_]�VJŅn�
�u�ꀀt5�+�ĉgy����l�-����9�n7 ��J��B����d��M[�2Hļ=>��R6\͉�����yz��6T8tX���YpΦ�e�a!u���~������f�E��&��(����>�������m�(e�V�[��U�6Q��3���I���,�v1�/+�Fj�Y�)���Dtmk���X��CBg�2����Cr^zF�<#���)��ǆy@���v��f6��a���Y��]x*UG��BՁ�Q�K���u��n�E8�u���Pȑ��9�J	y��r&��)���mIt��̚; ���0��&�=��QCw�&�R�G�{�^�z����Sߘ̌i���S�݄�@ ������-'~����պ�<��3�EdS��a��Sn�5C0���b�d<���/D��8�Ԗ��N9!�ilq!��7xŗ�3Jϭ�8Z�Rxz�|�R�����8�Kef����-��i7��`��Ӈ�1̬�=K�aS��j]L`��cW�Ws���\/>��/���&v�������#X�D�Zt�,a�x��/�\T�Ш���c<��^>����ĭjZ���|FL+^��Zϼ���9��(![.s9�����Vt�9��̧|��/ǐT��l��,�Y}�;EɈL���%O�E���W�=b�g�B8�L�4Dn
�-����i�8��X�ET��j^�/9��}���� Ȏ�o����!�t�,5��]4b�)T=�q���bR&�M�u/��;�v/Y������,b�@��eV����(w�����\�*f2ڑX��|я
`2'���Q���p�\G�"�>�����N���gP��ogK�I���̐�/p
�o���V���[�Z��������p�=8>��|�Tm�ܭܹ(���U�x�y�"�C��_+KGv&%��5���LcձNrP�[����4��̹'Q��+�����R͖��{x1}�`m_��R�;6�%
k�Y��> �e)�$3]��5\g��?��;ݗ��#�8$�{~&�Ɐ��6�
x&���J���R�\E��+v�,jv�\���s5�E�����6�=��a1D1?3][�/�r�ǳ�@ϼܠ��T ���/nֻ���:���J\��ȳ�f�V7�sB����w�����b���Ίz:x���m=�|�@%V01:�V���)��w�[����v�p��B^¬k�P����뢱:���1|Z�r���
0�3,oiv�ܭ���5�ij��j@��e��hP�r��"K>�.�}�a���+�����C��D���p�uOd`��H�Jd����Sr �$��še$��K., __��������� I�֋7�P,zq�C9�[?�N�u҆� 6L���aW�V$a�=����}׍A^N�*�
��XF��,n�'�^9��x��6�>[�Z���jQ2�٣��rt�!�g�Wq�l� ����F2p$rݻ�F*:���ܘi��|��)��ƆN��`g��%xh�w`�k���^�U4����s����fg��z���=�����&�:���͸	�8"c,����ތ��>FA����c{, ����f����u>��h������:�}��g�Z�;//���o4�-^i�(j�ā�7�m�W��r��Qc
����~ZehR_�;���=ߗ&����WrlX?o4���5#�㺭�hAΛL�|��SA��&�����i������y��1�Z{��.��X�ˢ�)��x`ٛ*ǙQ ~R��5I���ZŁ@��m}F����zLy�ؚ�,�)i��X�H�<��ťF5]�,�-r�&*?�z�<���S��q���9)��5AW�����i��3�1(�&�9�[t�M�{�fn�=qq�*,�CUx�2�9B�WJRSMȵ��䌩����E@*��T�Kv�%�/[����yr�Vz�c=E�������v`.�I��6r�<Ds�܎Ǹ�e�5�����
{6��M�x:2�e�������K滽G�1ip(�\!���`B��х���/���vo	��M!��ywĝ�Sf,v�[=����b�)��Q�I�p�V�@{��a�+����B_O��p�@�ϗ���?��FwZ��@-b�W�	j�d͑R����ܣ/`ח[����8p����	k�.ƒҙo�?53�͵&�]�.�b�tHj���xU��IQ	���ˬ������?Us�=/ �4��"�"K"��.���ש���q�Q�M�^b���2��������w�sx�S:�A.�\1x._��Cy���$�yT��lxIM�N�n:�?�&sG�?�q�X����������Jt4?g��eTQC0}��L��
�a����?���d
��5R�(y�2�D$��6�VVQ�>�O=s;��{�
%V�����#���������x	w�5�uW�s6��a�T������	�X�t�͗�-��{��mP�^xx��r���y�6I��P�L��j��n<\�� P���T>�����k�S���"�l{��ù��7)��ع�fx6׳9;`���m�W���l�>�d�e'k{Wu�-Q�-y"�a�Rn�3����F���"��:>9�
.5Ĵ[���<<UD�0�f�sCC�@R��>&��Xw�g2�;"���
�ܛ� ���*=�w؜�D�1� �Κ�:���I�,�E�|g�M{�#�0l%�/G������'K�7�A������)�u��!��z��Ԩ�Ҡ�w�$L#���D�3C�-r*�t{@�V� X��3���9'�	��������?V����.�� LJ�u��%>X��]�았f��L:��A���)a�[��\�%��bM�vv�D�W:R��*C�qM���?}�<#�?���*�[Kഖ�A����b�~08���vj�{�7�Ğ�v�9�a��7+��b0i[q��}nh
ǯ�����������~�>o�+�xC���T�k��O�G�>�!b^�|y���g��a|�c�����Q]�%ՠdJ{����Ս�1
e2�3�m�<��$E��E\~�����~�\Y�j�>���kM�'��oD�I0 ��z�P���|�ɞ�^�M�H�_���bwa�M��O�,�\&>�T!W�*�𥆐ܻa��殓��+,��;C�� �����d݌���ZC\9�/9�0Ҋ��
$v�(�u�������������B�w	��^E�K�ga$z�Q���?s��G��}������gee�|��2� <C ]���J"-� ��w���4��e"�5~�s���Z�C�>(;L���L �f�R�����T��+�Nr~����h����k���ڤT������P1�(:�3z��c���2���N����ɞD���R׹�کF�#����Q�4<�.�4%�{�����NS�\r�"6���R�=9�qh���R$4J:tb����iiv�c� +++uj�_�+3��9?���lw�߽�t]Q� ������Jco+���M͛'�=z�%<��\)5��:�?2�g4��,�e d@
�?2!U��iMU=cն���ưę��f�#R��i<��ZԘ���o-%��:G��*�z�D����p��>A~koO/;�ȓN
��^���
��lѱ'_5�Ճ�RZK�d`,�7�9WC0����Vp=�{���"Q�~q���:n�-��j�-R��|��c�0V��{i)Y��'
-'���I
�c/�$}
`F`<��s�.�/Ժ�|����奈���7R�[��.3���\����5h�;�,�}�J!�	6l�j�I��T�{�Wi�Ƨ���; �S���n'�қ!��E��yNz��F�\��E�c��ȹh[a|X�ޔo�*����.G�KҒJ%�������j��}������ H�^|�,ҥ$-↜ߧ��ʯ�;ie�/�th�uxܩ�a����8�e�'���sʻ�Ci��۶z��s�~!+�הּl����ysSKV�O���y�����$>���d2�`���I{�nL�m��y5/Tƅ���&�Ć�}�X<�e��~ߙ��GE�%������B��&|z�< �_g�'�2c	U����hvQ���}V
��D��x\l�Eb��
���X�-�m&�egw�����Wy�ǎP�`O����0�i�'�0s4 *�Q��w�n"o�f�øJ:%Q��+U�t�2�{V2x_Vo0�+��9-�[V�:�I��7�>�,�^��Յ9Nb�7�����Y;�U�u&p����b�lV��������{^_s-�Ջ�r΀C�٤�"��!+M*�-���y�$H�R��ʖ�F�W\�'��'׻-t9�M� ��b�!%����RI@ ����Aړ��] 8����UML2}{�)Eh�����3��m�����I�i����
 �{��X���A:�s'�~0O�j���Vh�Ӵ��ٱ��ra�/(���b W��#�3�%�xL=0R�����ׯ�N-4m@�ެI��D��N��ֹq�gl{��m����l=_��P����H��"�ܕ�]>Z��O����M�=�0�կ0��Dӑ���7���M�2}���O0��\i V��\r�ZL��i"���y7a]�<�ig�w��fN87P��E��==NtߖN�1Xu������P��ﴹ������x���#*��$�kÃ�蚮��e�F��}�3{�RQ��%BX1,�cJ{=�>..N�P��e4`�t�6ӭ/��� 3�+XZ1}���1 �ǩBZ�����Kä6���}�E����0:̤1����l [:�iD]~?��;���şt�b���f�;�<�]y�G*s+���Kȁ��˙c݋�i��Y���@J!:���W�҈��{N)0�������r|�X��Z��Z�B��J=�O �n��M��Sѱ��ԭ�7׀�8l=�8t?�0k2	D�S`��\���e�������$��/c��+�u+R!�W?����w+eO�t��
�+�
�����~�@W
����V��W�qݏBCt��~�@��6r	�@0��s��yb�M;!:����rE���PK   ���X�&�}[  y`  /   images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.png��W���x��,@���$$��[pw'h� xpww����]w���{��p�sf�L�tWwu�S�]���(�P@ ����2s��{����[�<�[��)Z���@tq&����醌����Q�ܕ�ã����0��Ќ�P"��b``�E��X����t��a9�檗�����EV�����*f7M�?!��ģ��JHH�`�s��m+�>=,?��8�B�ybѣo�h�I����7�.5.��}7�O�3�����1�]��fPz���	l5\B�zB���Ǡ�9�WQ���t��ԇ�t�D���=$9���y?����K=�`�?y.��d�bh�h�� ��;|4��e44Z7���A!Ɂ��Lс3N���R����BS����d�����_^��Fe�v�����t<����)^�"��y��(�N�Eİ �7�R���h@��`�(
��@�� Ё!ğ8��(	/�e$�A�]wb���?d)-g���#���(Dr�����C�G���!I�_��������{'{sK��.�f���P��z�>�7�Pz/x}�^�ʧ����f+%O)%�.V�>�9y 8�o�Y�ڢ�d4q}�o����V��؂g`�`࿘��u����_*�/M�ܛ�C�M��T��0=��������,�.^��_�������8&3E���1]����ߤaV*宣�K�W����?��P��|����������gi�j��fJeSk�$uQ��h�/ڳǠ��S���+M�x��}BM�9�+��rE�4dMӌ�����b�hp@���/fg�����Njy�|W"D��=P� �LC��˟@2b��+�U��=L;S[�1}?�	�c�'�z�ײn��Q��I�g���)�GD�!����3KWEc��Ǝ�YXG����w�W���qO�t���?�z,�����=#�Mp�����9Iq�����]fn�����\QQ8қU��X-�?�瞭���ܷ�Y�}x0���]���Y�c�����MY�W��Q����G�E\ж�aL��f�y(�3�_������ţ����6����)A�X�֕z�ΉJ+a��©�����\l���f:-��¹�/t ���'"�vy5��S��Y��u�èh�z��x�ۣ�ni{0xq�ʇ�|��_#[���%����*��5� ѬXX�'����K0y &�>�NTm��Q�׋E��j�@�	�����z�f7�*�������i�ǐ��	z�M��)+.���"}Ƙ�s��̥�b���93�R�R /�y5R��w�>�v������Fdt���v8���ډJ$J�ݜ��t�+�~�?<��la��綖Kц���x��+��0Z;H�fp�;����7.�c�sϋ����?L4j�ctҲՊB�뚚�&�n~��/H�X�A�uM�Y�����5�W���a奫�r��E��泑�'�'CR���:N^��#7�2�d&�o�ȩʓ��_���ne������;]V�	�%�R=r�G%N�UH	�|:��}�$�$SX9\:�H\�.)ah*-Ywkݸ��l7��TrCnElN9�����
��xwy�����=����$�a�V2?�I���)��5V��'<<'EI�I���%���-cO3:�u*b҈�Kl9�@V[�~%M���0`r�b$a�k�G�V����;-����m�'�{����6H��ca)��rw�p]�s'%���R�զ�ţ�L�L��Iծ���_�me$-:���y�'N|�ޔ /�B����(������\���y�I�f�f�~�ٸ�(ka��o�e�����{�)T�,K}!Q��`@6p���5A�`�҇��P_�3/A��8yZ,,,.1FF�Б}��'?�-_arFF��#��k\����~y�STf(JKI��efe�zQ<o��F8���>�!�lU�{�)�p�w���,.vj|?�!܉)_�1���ϼ��+{HQ�W�gmq��@WB�`aVN�)A,��<�:�^�Y��CJ,޸��o(ǜ ů��gwm�@���8Xt:U�.�3/_V�X@Bs���8�&�3�`^?�k�of�Z�0���%��2IL�P�������d�*�5�-M=���m�D��I@�)4�
�wQv".#(t"���k���R��,�WR�	 �ϓGEe%P=|��^;��_I+[kRk����J~��(�:I ����|8��d��%���z2=1�+�u���k!�p�P/>�/#�e�4�������5��D��t��*ɟ���8L�WD0�OD�(ɀ�6�a]V*�,_�r�קbC4�\ $�1�xJ,SR�r��z���oTgdS�[���C���m�:-���5�t��I
�KͿBʜ^%�*��'�����4f���Q(`���u
hR\.
���쳜��dMV�#�������IW=��x��1�ʐ�ߢ��3�����B�%L�D��!4�0+M��f�3���o��&x��-����Tl��d2��%E��`W걆���	�ε�O}�!9b��7���ʷ5���$˛j.�����K�8�j����#�psJ�{"��<|��[�v̆[�mIR+�?v��psL"��kDs�X��ݕ���)����2�_0E���c�3��Ȫ���ϧ����t;�	
�UUUlbb���n�F
66,�jA���IL]N���ē�E���((s�ak,)d o�~��oR��}�Ku=<��1��Y��t����K;y�V"(���n>��0��W+���,�P���sB.+ܚv�iND7J�M����w�r3����'{
���k�����-���4�j�cm\|\Ѿ�o�s(��+�cz;�7�������ⶳGԡ�5̙�~����@8�.c��m�� XE]m��� �0��a>�7}eY�՛ł'�äa�.<�L��ۄNm}.���0s������O�TUL��#�\�������.'z�	�:ڽa����H���x:N���w�ng�4���$�S����',x@���2m�]ەt�QO�ϧ��zkZ������ HS�f���`�eg_�;��l&F�� ��۪�� 0�A~�����{8ܙ%I�[��������灚��|��<��':�N��o��P�4L�Q�z�������4�c.�{6�?�2 ��U�Tv_�&y��v�G	?����W���4�apP;A��U�4�K$�ԧBG7�%[��r�6k�n4l4��i����=���d�0�����V���`���C��s)I�=�%/�4�u�9H���Q����'�,W��ЮY�B^ī܀��;��@��T烌(�7���v���98��Zݾ��1�����78HEC�xR�����J��	E'��=����Ϫ@*�^/+�:*��-�C������r�(�*�~3鄖>{�q�/���f�H�ܐyV]/�����ްd7��r�ߦ��0 �jfjn<:_���2CYV��Ç]V�v��+t��%s��k
/�w�{&[�s\4�)A�k�=�v���-7�#7DW�������"��yZ �2n����Ir_�ʗC��62B�̘�<�t~_�����Q�l$Ȏ����%>�=v��TpZDD���M�Y-�IF�/�pq�{Y���<���s�OW��Ef��iΉN���ߥH�:�0���(�8�n�5;�����;w�+�O�e:OG����\{�B��S��h8B�ޅK��NC?:=\K�{�����x�?#U9l|^}��r��'��c��)�=�Y��F"�쩅��h�n�x�ﱿ���ܼ��B��˧�pPx�����C�!��Gx��|�%���5Uq���pH��}*��^�{V��cq៞=����U>9��e�~�	��b�u2�++��pR�ȼ�굺�9J�ޞZdn��w��g�C����R�sB�x)�vb��/WS�֘Em?`�r,���]�<��C��H%�>�b��)�13tɰt�?}�2���x��iz��V;R}�s���7���&g?)�]�>^�>����c�����X6������I~�I�%���5EA�N���l�b���ͪ�\�N+>kr� 77���H=!��<���,�-0ߕ��D��II���"aK[|�|�3�e�_��z�;�hO���a[~���`�Lb��e6#H����M�M���*Hd��.^�$`�8�{=�r�w��K�~�y�b�x��>o\>l�{m�`/�y-w)�z)�ym����8I��N����[ �:x/�=<Ui~��.��*gM�E�77��El?x��{�&&nظ`X�iؠi��n_ن�8�p���n�t�Ab��K�Pd\;����.��o���BU� Y�%F��Bp&>�ß���]����k�k����ֵ�}�APy����5���K�M�K��k���r��jIy(C��EO��N�/��+��sU���ؔ�¸������Z�x�<A��u����d��:����t�`����zC�W��_e�.���������vY�S23cA�r����(hi�ظu��뒦/�T�չ�Z�M?ub�F�(n�f�-�u��>��f'L�������0��:����d����!�J"F����g��ɜǒ��9�*�a�2�F���������d||��>��hd����T��cw��J?~\�ή�Y��no�j2���dd`�n�>R~mH��D�ݦo�>?0�#�����c��E�jR��� X��<xkpE�fd��
��b=*�2 a�SW'@#��E�������|m��R~L.D��8��\��ݿ�Zj����'����ic�����'�B�5�% ����0���[�΅ʒ��Җ�3�I�R�R�_����)8��LLK�\����o�!�����~���x���C���?	E#z~��*�f�.ɫÕO*�q��ɡ�]4�+)j�n	�ܪ;/������g1e�I��Ӣ	@����n���v���}f!S��G,��"�\V�[��X�|
fa��"�L#K(i�X���|��S���r���^������G��R(���O���moMR��t�Z�8n>����U�!¯﹣�v7��76I���x�y_�B�������n���>?��|	J�+č��YSF!��8�|(��|f�C�V��d>�{�U�w(�xx�
�ď*�i��=Ճ���,��1B7�}|$������8%�A�G���j?�KȥBIy^���m�7�-.�(���EA3��3Ӭ��ot���m���Ә�N'&�2��ڣ�e~ge�'oY��/%���$t��j:�Y3ꉠ}�F��殺!��`��xg����ua6���T���w��j�2��KX�Rh8��2Yn�F�Ie8y��2_�&/))�R]�N,��M� *�� ���v{68?i=5�nD�2��ed�:�'3�h#"ƻpz�Bと}�R!&�����'4��[�oڮMJ�����������b��$?�_X�78���؋�U�D*�H$ǁ���I_�Dz�ɳ������]\\�L�z�����̒,eL�s���ꏈ�^K�G�L�?��.��a����贼�6��z�"��\�ęq^�_�*��q�h��{�c{����y�
q/mw���0��2w*�`��Ĕ�/ Q�4�����;M[
��L!X���kt��k��
�,	������D�qh�?4���r1�U<��֘썫�M��d�q`�+o�����4�3'^��S��$�vUGGG&9���Ե�`����_B`�����
�V��@C=��d@A�mk=�:i�ޙ���A%�oe���^�c��~_T}q$�B���".�g�de{��qX���.�􎏅{(~�<����r��ŢǴ�?L	��7��C�fo/,c��R���&kπw�o�ӿM[P߾Ϥ/���宥34N#�Me�O����l���O�MFe��z�Aڊ�G���p\H$��g ��4��[&�D���5)=�gRS3��}�
�f�fn�V�����T������bꞘX�.�g���^�����$2G;���M���
��`JJj3����2{QeU?�rS���fL�Z\�����tfV5��	�wk
"s�I��Ѳ#n2�_S&c;?0��{�6�}(��r�KZ���H�|;��& �����kdw�6��>�tC��-Kwк��R��˵���v�VzWhi�џ$^҉�	�:��l�s��am�ߞ��Cn4�	!�J]�����X�'Zī_��>�a�����zQª¸9�����B/n�Y^��.>��������4��� JBq���P9�W��+���'$�J�Z�T�L=�J�2B��B�x[7��_��/v�aTv~�K|闦k�g2��W���Z���صh�T�{m���:ָ=�/��W�%x�dP#G�d��(��4�K[�%���}�W�Tg.��� ��|<m�����P����"�y�9BIy1�s�g�Hv�v];,��n[���D��7X���?vi3��b��A����>_��9�ȸP�#�:8ty������/�+:�g^�~e'k�ħ"v���Z�����Z��{j�#���_���
�d�wJ�Q���N;�F*��*`S�"&��V����{�y��V�Hs�y�b�8\��~/7V���o*�֎j6v#g�{�#,�E�,��-��d�K7
�8nFA(�k�]%��TA������	����E�ʭ���Z��ʦi�D}/df��vB0RǮa�qw.�rx�pZݹbp`��<�Xx���I@�"W���b0;}�n��ZA䅤q���fM���~"onb�p�K���a��#����V�Ksj��l�Y�W�cBw���!ʋ6�\���3[��������|�}�ƃ[+)zP��,�UC�R�?9ϲ��=�g9�Rμ�|���@B>'ܚ�������EM��У���*���Gk��-�U��7��MwiF�K�����*,��ka` p\��;ط#n3�^�̗����D3/�%'�e����&�*�&�v=TWm��`���<_f�����֣L���fH*]u�%���tj��ҨԗRP����e&p;��p=A+V�2z�&��56���cf&xI��C�%?c�A�<N3�7�ԸEHij�R +��@s�)(`����,q.lؚ�E�*�۠��[����A@�����s;Rh ����d�x�g-mup��o��h�N8󜳿e-��~�pvlv�JL��aI�~��+aӿ(	3O�I�!3�,Q����#Qp1�;VW;4��}�(��O�Ϭ�z�/�,/O�|�i��%,���h��ƐF��>N��@8�C� �@+* #�\ ��sz�%����Ca?�����]���Ȫl�0�
M6�P��uϐRn�e�A'�W��B����څ�U� >�,䝚ʕ�=�	P�yO(h:?�]�\�@��zb����Se@Iy�y��yh%��SR���_:I=�(kl�Q���\8Ԅ~^�g씈�Q�v��_����AeL ���i|��d�c��ijfƣ"��/b���j�������(���{��q���Vl����FiG�&!��{��s���en�Տ)T���hZ;f�Z���ӵ�w��
	3�"*��l���22��)̫S�gѣi\s,��vAM��U#�r+r�,cT[e5�5��"��&����js)��ǓQk�Ro���h�6�>d�{d��T9�b�˒uڔ�1[���Qr��y�t|��e�3�5��l.����kA�޷{A�}W��}m7��}�;_�î�1PcE��.�k\0��Z�	+'h[�'��"w��O�^��3�#b&�t֗�Ǆ;&�*�H��'�]���i������K�C����umm'M �\�M�3.�%�G��2XΑ������H虙�d;`�[�Gq+�п'B�fk�p ,[�u��~PU�ɩ�ڍTc���eq�ys��9=n@����`�S� ��-ڎ͞�s|��9�)o�` 3X������ܺnG���;��RJ���ݧ��8���[;���+t�[�SR��)�������%w���ݜ,�=��@�����3�j���-�x��6�.8��4ᤎ%,�4f�=��30[�	�g*<?�����ɱ���UDw�Ɔ龠f��Rѹ!�Pg&�hg�����xFg���V75"�Y>�->���Ѧ\�ݑp�\�������Et�R�h"���:���3E�͑�ne��c�g���4�Au���˼,��-zc��429��/1"FA>���JX�����iX�n�]��g�����E�I�w����#"�?�yYY���t�H��u�K���sz@J����=�{Mm%~���lg��I��5݆�%Ɗ�0�3��FcI��1�`Y����Z����2��b��y'~;G�4I��[��eU������׎Z�G�*V\e�zM�s����^�!T�Y?��c����_q_���Z�) ��村���!?���w<���S��t��G�9�rc0s�$�5a�彐��|̯���?�vC������m�<��6v(��ZҐ�:��~K�����>�i�+�Ҿ"E!�$��Q��A���r�|����Ö��:��7��K�����Ճ�P�eWa?׽�u���Sޜ���bL����I�ZUL�y����\��e�۹�"�p��`���x�l�'�K�}!���Na�� x��Sn׋j����BQa�y��V��1_tbn;�A�l��z�����T�zM��0����¾^�2��B/M�8��7��f���n�h�m�tC��c:�L�.��͒��5�',���/w��}���%́�����MO�Kl&�œڬ� ���s���K��\Ee� �������+�k�RU1�A}y��~��M�O��:.h֡^l�!�����[���s}��/�Znv�vWܐ>�Z&{��.����)m�!���_��:�S+j���>���f*ii-<V�(Z�L>n$u�h`��5�A�GD1s�����z5�o��!C�����n��7'+�D0�\č�~�����$"tkpE���:�l��#e�w�p�is?��i(��a�?��8�%$З�%n���"�ܔ��Š�\Re&��Bj2�?���['2�\z��o_������P��t�}���#0�m����J}�"�_���c*ӦF���s�t�ڎ�=�.Ǳq1��KM`��j'��9�"��]E�J�迬��a���3[�ˆ���%�U8��|.B�
j�F폼�e��zk�(;����쪢"=e��BK�F�k)�������_	\c���B3�/·�bM�x��5mo{�_�b��KK�$��\�zHaT��& �P���9����Y�@�kZEE�	CT]?����u� �c"����������I�#`�U�Gd�R:םqm�z*�(��H��QaM�ڮ��2�r� �I>��;\����aGo��cf�d������l��t�k����!m�]3@���mM?U�DH��BF� 	7�wqOD���@�:�w1?��g<��;��%�㚰/�)D�*�#RI_�Fq�?lQN��T���,F�p%A�.l�
�~^á��j���gɵ_�q>���b�%8؝���@,*�H�
W���]]b�����3���Z�	=EK�"��9xk����ۖ�����r?�AYI	K]�3�g5W�F��Z�ZZ��gypE#��(!��=}(���gX~��&�/_�.)�N;ol�ޖ�رk9<��Q��4���N�	��Z���t>5��|�m�W�b!�`.g=3V
���3�z�c�_۽͈K�Zbw��2h�u�4�P��,�V�m��h����t�+]Б�K���� ��T3�|�_��������ݞ�> �$��3qm��-�p�~ 0���E8m%&/�C/4�uM�g��5ب7��=�ưZ�g\�Q��iV�٢E�im1
��NN_�}{��!��t�gy��j[5����v�E�X�ڲ���#��LH�*�zw�Iҕ����������$\�h�5Pn֔����%�E�ʢ~q��k�>ߒӠr/�	Cq�x�m�俙t�q>��M.�r���eu��LS�v/A\>j������2X&�����,{0dOy�#�oY��UJJ��-���q�{�F��CۤE�|YB�o����:�g8����������!�Y�>���c޺����_p0�0�B�0�� �H_.q�-��NP�qɾ��c�-��wD
6���.e����m�R"9aa�0�����IP�ԗB�|`�1��(��ZD�v�ߚ*�Z\>u�=ah�kq?]��'��=��&��Ňg�@�>Zح�JEl�,��@KK�*��h2�s�����eU��~�o{��e��ȭ������T��w�����qTjR#�7�$P	�b��{�dLwU��IS�ݵ:K�4{�D�l��?U�K��l���g��A1�a�D�RK�N�369��d��#9g,OΔ55�3�	;�j5�vmPa~����!���e�-�~l5���D �>6�r i��i���wY>y���ɍ�$��4S6�V�3i�&/I~��AT�_o=5�����1s��]����<��\�F;֖�V��ӵ��v��#7Ss����ZͲ����<Q��5XRUc���pRah�����T� ��KVI�]���'Y����U��+--r~�;t�}��' ΐ]ˊּ��f:���vQ�GWpskc�l֑���������h���/��$LH�C=� }a����Vg�⟕";��N�����J�z��UF&;{�DQY7�'���vЪ����YoƎ;%���[/���j�{\>}��¤�y�M`Ż�]<�"��**��03��ʚs �9ɕ����~�����(~��H7�LYƤ�a���G7ɽV>A���-��56U�K�Y�;��O~$�����d��c��y�'��0)�5�������z\jHr2%K���&?Q��wؽ��%�.�cN���~��s�ϐB�¹sPRWW_)�?�C�M-�z�����TGm��^욐�X�aŭc�F�(Z��O}xc�9����7h�Է��(���F�%��{y�����I�3߰��+l��]��Xܰ�+F���)����)`�Q�<hI��������Ia�S(�D6�c}Jl���O�I^�����1e��y�G?\]_��D�Tx�v�ȫ�Vѐq��>�N���C���mv�y��q�-���Y\BteU���^�=�L�{8�h|A����[�W�ݾ1����)H���r�m�NVr>%��Q�Chu�K�'�7�h~ˆ$�I��e���l���SD	I�Zs[Օ��ދDF%U]4=p/���	!yj�T�_��N��X���V5d�;��k2&	=<F��!����e\���>����z�$B�s&yL���P�$d�o"�K��%�-��D�a���p4�����''6�[�(>�W� /����m��7�_@��o V�R��>��Խ�,�2�9obleQEiU>)����qu�"0)�<��hΞ-�Č5N����V�Y�-ɟ��"&qtt,��|=���X�����-,�{1�����N�A�5��I�|���n]ƇD3;|Y��ޤ��Kᵚ-�ӷ�!�[���y��ɡ,s��	$m+QR)���i`K� c�:E�l�yuU�g���s��C:���R�3�=m!�r����ҥ�oS=�H. �N?�����_�%C��.�|u�:t�H����JD[],����r�z}�J��m{\�ޗ����lU,�m�h� �b)
���h�ؒ���L`lB
���W[GS.Δ�vB���m�<�����|v^��w�R�����֮۝��Yb+ ꀭ������*+SAN��Gb���z����f�V�M� v|�����*sj�Ȅ#mLJ�'�_>;/�KH���� ��_��:p�v� �R�xZ��6��Q�kL�f#I�3P�l���3?�qDޞAVJ5&�g�5b�����Bщ�]����c�aׇ�>��G��%���#	��Y���r�S)-kCp?�ra�ЖE�w5!u����C��y�C��|�5��71Ye#��=y��90�]��rk<:6��d�޼�QQQ��0̖Z��D�`�dH ߛ`<�;:򁚺a��H�]�j�W�ym�>zY��~�}$A��%�\�c�tDMj�\�*�oX��2f=V��tcE�ҘW��d�u�LF	,9�Y�@%SP��!ί�� �=��A��QP���[(�v��p|���R�m/��XN�")��`�+KN�j� <O�'�G�?�SSS?�Vh�6�j6#4�-��l7���C����hpQ��L��L����:�#��;�W�<�&x1��������ؘ��b<����3��z�zu�4Xe;n�m�Q�Ҵ�Ԩ����q���g��lN���t������1<����s��v3޵��-r���5�1���U/���D�D�!�,͸<˷��ɳݶF%Uվ.y&ʀoo����_1�ð~[M�����z�6���A��C�J���w7�ᱳ��~I�=���D�����!a���`�X�eP��Ю���z��tp���ſ��m�@��lQ�t��w���tw2���G͍��d{���p�H���5�H_o��uI��������~��qd�g�Z�\��N79�b���?��Qӌ1���ɔj�Z��2/�I�:�B�VE`
#���Ȯ��芰���]����b����Xma�U�گ	��~���e��	s�%�9�=��^�LT���}{5v	@kҾ弘�<K��<d)i�w�Z��~��2�떠�0EE.�k/�<(�Y'���2&1���w���eip8��k~�uz�DЌ����q��6���7�{X�5w��������=�`7+��"�;�K�F�;(�����!�׌�|/O��G��KR����-{�$�A����n/sɬ7 �T}��0S���,�;��h��rhx\x����[4J�D�糀
��R����j��g��k���F|��.�02��M����7���X�!��(˟_!m*������V���[��7����EN��0�}F��ӓ�v�z���vm/S�M�
`é��P����̯G�X�MfU}�苠�0���\�\~y�`k=#H�y��P�\�:��\aL�J��@�~�jȢ�\���^&��I��/ (�E.~���/����g���EU �z��A��\�(o�Ջe�iLo~C�bi�qq���d�f�H�E���Z�_~.U�!	�&���e>�2�@�_ױ�~��t�_au�	.�BE�N_��e�P���ey�;�6���|���8��'�`c�j�v����3�m��\�[e%[v:�D�M�5~8���X��~:�˙�ͦ�ذ��k���ډ��0��J����^�k�{���J{j�>�3w>:�|�9|��]F�ϭSE�'H��Ϥ;18Ȕ���o���X�ҹ�J��j��[�i�1�F�;31?��x��Gj��	qM����> ��v<8ތ:�A�b);��xq���ص/�5_*��>��&�����A�r1����[X4A���SV7ç�-�ȳ�Ê�N��6�������0F�N���'���Y*��*ZOX�F���7��Ⱥ�xV�����XK��xK]�{��z3+�P���{���Иl��Se0������!�� ��h�z��^x��4:�Iؠ�W��F������K��T/]��^��;.�i��}�"�'+�[E�1=UbS���ff�DF����IO�WUW7~y�լ6��͢�/�d��`;�[��Ubu[��]����JF~oII��D��[��w~�}���$~6�a`�������p����Ȃ��TP�3��s6Fntb]it��mѕ+?W'�O�q��d�w#��v�P��fD��5��V���U�jQ��Fb�Awe�����ȉ5��aY���Ԗ�x�\�M���,7Ϸ9���B]�O_�1�I�)������/���)��B-��������q���ME���~~0��D7�U��b ��gs{n_a�0���7u������-�%��t�ѳ��~�Qe��e��Df�aڻ!j��M��t�M�դ�̛!����[SS��XaTc��6�95H�]�E��;
���ȡ��e�����'�W��ĉ�����.�= m6^80G\\x4rbFJX7�Ka��2��?�lB��g�;�����CF2��f6o�l 2��?������O��C��ͷ�,��R�͘%��t>g �9��W%�����-~8����h��Q��Ͼ���_��:����iz\��i�$�)+X�-9y؉��z!��E�jV��$y[l��-���S3�`�%�wU�Ԯɂ�a{�!X��oap�9��t�T�]���`מd�$2��v�0���聕��b~�`��c�P�k	C�̤.+p���}*D(�`ؚ��R(z��0��h���O�����gE��*�s�_�z�Q�I�k��9bh�း�������y+*s��̭Y�wyP��S�N�J�����r�޵�4�,�3�qo�����Y��d�C���Z{۰�S|��+��ilT�4�)�o��m�>�sa
���{����d����M꤬��N��{��\7�g� }ot?Z;��X�53!wC��4G\�<߭��,��~KԴ��v��<Q�Ê��au��J�斈*�^�v�J�\	F�0�f`d�8��=e�a:{��E!v>����p��)�G��ѡ�'��ÊF��_X�޺�¨�v�@e T�)a�p]���	�!�ޘ�$�N���(ퟦ��J��wW�a=s�pQ..�_��hE�m$M
l��w���m��e�(Vo��S:�"��A�}KR��~��vq��t9.�31n�Dg&��X�p=Qà�����9r�щF�d3�IJ�k�Y�A�����'�G�!"��$�UX+��_����0-���:9�!ÙuQ.(�̺O��Q������t�UϪ�r�հ�a�7���/��d�4�>i��Ɛƭ�|ñ#��r�-��|<��ܦ�?_�>��]\�V�U�֎�+o�7��Џl&돨����V��|��R 4R�7���
��mA_P	�k���'��ǒ�N(1B'��.S!ɜ��؛����v��.��{�@�של�o�ݬJ�����'���%-�<k>DvAz��ZW������Emdј�����_7s�}�`.��O`��D��=g���0^����enZ�1T��RO|�R�������O�-����w��Z�^^���h $��P�`�0�#�`u�F~��>�)XIq���ѳ�W�\�Ez=9���}�Y�D��p��x����P����
�4b�z�Ί��><,�k%�xW(ˏ�+#n��= ��y�
{�N�|�}m�vBx0�j��3/��:���hxt�X�~;�	�&3�>s�_��7wh*(|��5��r\;c��;XS���YU���۠���Ki�HA��Ֆ�A�h�d,�
�Ǚⷂ����voW��""Bn�xbg=p\Z��
�[JJ
!��G|�aK���}�Uu�qy4]Hz_��x�TC!Y[oD�j.j�l���qz�Opy>^3�>P�b	X:�p����cll�JO��U\(ߋLKx��<մ���S4rn4555tfePB�*/��z���I(я��_�k,X��[?&ϗ�q��&a̫�ZM��w��P7��d�Օq�Ё��Ns�����;+�'��s�kk�OWjgϲ�������^Ū��9��T_�^k����jB�����p�<���[��܌a��ϟo_S5M-,�xx^��gZ	�g�+��\?Zݔ�=�!��{�/�oG�i��~B0&bc+J@�uu?�spL՟�w�׻�����C��~o��@���:��������u�j���Cs����#ŔC�AT~gg'��[+���y(��ƾKNM%�ۼ�HZZ:�ס���3:>[��ׯ6I�	II�;N�,gO�o^O���ޜV�Y�A8W.�VY�+�ܛj���R(������deŁ���p]��dU��]�G�$�F`�t��p�Bs�����k�7��J���\t��q��q�j�C�(k�E��m��3Z^���ˋ��R��!e�%�!hi�n-�y��Ã^x�f�U�p�И�ZB��QE���5�p ��bs��b������w�!x���z�� �db�0|���,���u��D�E�4ld'hi+���k������������mfq���:,�o�^��3��
<"s�yX����/1 ��ǐ�[��y5�P��*��bM��!�XF���9�����
*��Z8��Fip6�6�5��tMm���h��!͵e �G��|��e�!�]�)!�{�E�з�8Yi#fo_�l-�.���~6��G���z#� b�ye�DDN��_�{���_��>�8�zK�,�_��FH�����ɇ\���gV�|EG��<�1���Q	)��H�������v�ɿL�T����e���
���OG�TF*>?�g����=�u�^�+g�{��#����Ys^iRÈ��B����K�Ķ4��BeO}�4�a���y���n,��S����_!Q��
J����B���K:M�f�����]}V� �����.���kk�qg�͵�O;���D����
�4�]A@ HP�Hҫ� RC��(�{G�A��A�� -t��J w�����s����ݜ���}�=�<3����Бk��Ln�Zp=�.旐�/9�oڟ���ƶV����"���2�=��$ߧrNq�9���2w�|w��ר����T��&Ӷ��MR�G7g�{,���gl��W1�X���_%z�"�����-9�`����_^ِkf��;/�s���9B�^i2�,��&�m.��hN
y��2��ry��/��ƫb�L�����o�V.��ug5�"��x�y�m��N��'�)�)���-������az�H��}��Q�Ļr���3Z��̱�g0{��	��*�V�/�u*v�����1�|{�l1��.j�ɠ�.�[�1E��æ���(���$-����=ط����k,4i�||`��3Qi��s����師��B�S�Er&Q��d}rN��	���f@�g���@)[=�?�2�ݿ�&*���+�}��Y\\,"*��j-q��n�%&Ջt`-^��o��W ���7V��ƪ������۾�HZLѰ����B����QO����Se2��><�����h����&���������S��ތ5��Q��P���-�LHi�Q�]ޗ�WA&�3Q��Hr�U([+��<մeҷ����$;�k���X�ys�a�� �b�c�.-�Lh~tݟ�t��)y����]ccc7��c��5������F�P[����~T,k�:�mu�t������[y�|�O�l���]�*�/�b�$�(��Oi�`���q��'^�e��D�-��$�q���Qjt;����`�	�G�؇���s��8H�3aTI?q����`�39�����RBɝ�L�������x��l)���*k�V���ې�O�W��L�e��8�s�K�ɫ���@�S���-(���ȃ�h���O�e$ě%?u�1a��Sv�m�cwĚ��La��X�ZkV���s�p��T��93�::����w���'�m�ȴ�4�������kWW�t���t��'~k#��=��l�cv5���ו��MT���"Sp
QśUo���a��'1�O�=����{Qk���
����7��Y�zEE�~�7a��B�aޑ![gG̈́~Y\���pe,�d��w=F�+m9�l�Oj�3����4X�mxL9�	c�������r�^
��_
���.'�Z��8��������C]{�1�<���7�D������)�Ϋw4����d�,�f�/���씙���H�Iv:.����˟��Lyeanp�⹫���y��+���1�	��je�\}�bO]����g+��Q�Q������5u��b��d��=ςPp+|=v�;S�C9U}��TX�5ex�*kc�~S6Y������W}=��ӭ.eZ���&y�sx�0r���L:�/�(H��U�^+�-�t�h�Vii�?4��(K��>c��(W�����8�ZA:eE����-*.E���3�[�M�z�uk6��d=5��]w��xP{������|�P(�w�t��5twT@�����M9��n���&cuF���ju�Y��0�k�rnM���S>!-��;DF�.˺n��ڻ{�;�5�#����{�u'���S�j�����t"A)L�;��G@�t` ���hű��o���b)��Z��jas�����R�<���5Nt]M�c�y?N���d��2��a+��Ɉ�)�|+��)���ͩ��.���\��lD�Z�[�����'Jy�o�Ve�[[�U}Bm.ȮU��g�^�3�)�f�׈��,����������!�x��ֵ�Ͼ���1��l���P��lױ;>�٩@O�˯'/'.�S7s;%U��1�P��^��c�vD�񭣘��C�˃M�������]�k�,u�o
;aC.J��~<���zÕ���������h� .���(��,ش(zU;`�3J�ZI�U���e�ƴ���{�Q�ՐLk|+A{�C���k��h$=��p������@5��{�p�U�1Z^_�'����KH�k�^teY\�u��P���i�+��g�h�^G���UCT�J��/�k��y)��6�E�'<R�za	��������]T�|Rq�����1o�֑Z��Z��-���%e[)p��#"(����JJ�`�7�u����8F��hx�}{�Z��)9^�"}h�6>�$!+mo�Y8g��l9'&6��\�o,�H��6f�,<ג2S��=�7��!(��������b�T4t�p���޿�O�+y��gf�SU�2U)-�!�NҾF-%�{��2���w����U ��*��H���Zt�|o__�f�'�`ȳݰ�^�������ԴTۣR�m5#7���z�0c��E�8׳�5�ظB~���z\�b!�c�֙a�l�ܖu-6duoxh��d������}G�=7�5E���qs�=ѽ����$7���K������)��/1�,3{e���+�,IIIrb#�m�'%�������i���ui�[;/�Bo����`���ǿ�"�&��f�}��
V��]Z�^8��9|.�sĘ�ƾ�q������m��r��˨��g3���O�v�gEEE��KŚɥ��7=>�W��-J�Fvp<���4q��m�e�\�<:�����A����M>>��s?r���g�E������k��u���Wűz��L�����(��:vj�j��f}@ژ�ԝ�^�E��	:�כ�%&}��!�UUؒ-�ћz���������	�E�O���y�2�F�W�����~ȶؤK]437	����܉�8ڙa�a��p&RD������s«��r�e��1�e������	���Q�<�f*�^�$�S��RRپ>>\����/�/��T�j��+!�|�"����#*-(t�ǚ'��#L#�kx��ƒzx��E�l���z�o�"t�L0��x�gD�&�X#"�jVPPд%$�(�������r��֝�bQAal���/���B�_�6��YT�� ���@��+��
%�1Xz�Cj<׎�Q��R�1� I�e˼�F#�<F�Tvo��f�ƅ_��|���2�-�[C���:E�ׁ����{e�+'��-!�Zl����u���>D�3���P���>]/ 8?�u��7zЇBB��s)�*-!v����i�^:���MuJ{Y���]�"�����x~�4�Т��R'�R~9� ���{Ff�ERR��������?�l�I~}�޼��4�B�*9[�0V�z�U�/�<'�\~���,�R
V.N�|���W�R���ba$S.�|����S�._߲�ކ�s]3��w'+�+�����<h-�4��|��.��gW'��q�7�s�?�p�|4���]��*���2Շ�_K�f��Z���z��h�s뱝ݻ#B�㹕p���l��������1Ny/0G�Z�Nf-�+I��sj,��¥Ug�d�J�l?G�.����,?�wEi)PD�I��ܹ
��mw�v|Qt�y���s7/��0��}���N��«V���弪L\�nf.������o8�Ǔ3Sw�ϫaO������W���mgvTU{���vJ��/���Q�S�Ҫ�2��-_3W[�b����w��V���hu�x�hXr?5"�8pg.��[���e y*������\1�/�4��k%�/#��⾩��}��GĹ�L"��><�]������+��e� �i@
���:���b*��ꇨ���Gbn���(�A6Y��i|�bv���u����A\כ�����*&E���+�q�o��?��r�70h�K<Zl"�GW�KQ�oQ�:C��*Vڟ�1�l{ܰK�.�?#p1ƽɜt>�~�Х��N�&�m�ƮYK�c9'�}a�x�k�A�^'�����~�������.������*Hdff6��qRڇ�y��֛�`�	::��i�Z��m]���X��j����5��0k	��h��L�S�+3�K���n^`��L�7�t���A%l@k�k��V�n��OgZmA�C���l�Z�(�����ȕ�yߕ���α����C>��|����Ze���9�Sq�(��˩���k��P�R^����n��p�@Ս5���KUؙ���>9M���[[�����+@�I_�����w����0\�s��HW������G��G���kp� �'�ؿM^�h������H ����uʝkq�{"�56��$:KMW	]����!a�Ȇ��_G9,�������b�A��X-��=]]k����t���x{ץk�G�a�M�;��G���U�HO�����fC!���C3iǅ���xxy�^���m�A��ee�4M���Ȟ�nd4�m@~eP>h&���t���{K4��>�/t(?��ܽ>H�Lܛ�{}�`�Lf��뛎�<)lt���n��I���z\ߘn&R� ��ܡQ���{�@�b �|��÷�Rls��V]�����f4���
��T	���*���*vZJ��xLCN+|���o)�91��62� űKo�c�K8����W�����F�a�A�m�Ɇ[R�4�(휗+}2� �*��M^+��n9<˯��Vڗq�%_��y�uq݈K/F k�D�C֋����}%�xȒ���o���eGgqX��B���W����y��Oţ/�Z�g �އl��K@�&Ox������xT^ʗ+8^��������s��zc���X6�%���P�Z�	��Ǘ�\����@H?��g��\H��\��s���L������_by�����g��t-1R(Y����R�4�m�y;��8���㸼�V�����r=�v��TO)=���6�X��\��*x8���n�cd{�۸�O����9S�4��@!7H�MG����i>{�\vM���]���u�ܶ9�5E��jk{{��JN���Ae��)�fq�Z�x��[B	le���۸�IN=�+V��x!�CA�*ЦJ�w�{�6�s�w7�-��ͬ|�%	�VLMq��4�(j��U�1�95;�ۈtť��+C��E�'���/7���Y�y%�Z3n�c���:��
9���ٳ�T�j�q�h����}���r�ͣ�!1��d�����Z���8�?���%�4All[���
�=6�����W�8�}<��4��Y�φ��s�;2�یL򳒲��P���ɺi�_�.�3&~�g���>���4a�	��_΍�\����<�'%%e6ό07��ݽ1]8Z�O�T�`V��ds��Ƿ/�)����/(Z#�e�	�x1�����c�N��r�Of� vP&�&Y���r-�_y�Ʊ؄	*X5Fڰ���|D�$O?�΄0��b+%%�����R]Ĵ]�3�h�ƈU��I0#��{ǘ+������݄���o�Ĕ��l��M"i����ʼ�X����n��:H!(��|׸�B�a�Uj����&����N����[����AK4�\�f�_�#����S����;|��w)���+5�;2�<)��Zj�>����\8�F���������KVψ�
�N�*!]f��g�V8L��Vm�z�&�$N��Qg�-�A	)9���dN�Q�-�>	��S��g^�/[�r�sȋ���8��l7)�!�^|��� [��$�y.�CU�~��}�V|�Q@��!��xГ*�|g�ۂy�ש�~6daA�H(;ؕ3��W�Yf��+7;y.,�Ը82�S�>�z#_0ao���'�N�V�?PXd�&�S�;x9��i����m����m�HI��}�Q�_JI9@�+[��/bS鱕���O�KY�|0|n���W:�]ٵ&<L�����[#E-��3��ɋ��J�s�"�Bl�GӍ�_�����>�)�=��� �Ƙ����r�k�#Oó�KVX�B��.����>��I	�����X NQ����b
����
���ι�g��'��pn�.E��,���u�����-�ԍ6�]ʲ͆��/���Tn7ݑ�w�t�L����r_&������Sz4SR�ϟ��;:~����B����GS��S�z��?��oI4�m-�QLwA P�������*>��`Q���~ 
v��0�E��0�B�J(:��}󿛬����{�,��W�ڳ���0Y���p�������>��	tC򆤸����ԃR`i)���5II���AOP���������D������E 9�c �	���99�:�A
�f/����l�y�tt7U�=r���yz�����9ہ��X�����KJ~_�JdD�20{{���W�����o�玗��#������I)9�6� ���8���>0/89IU����� }����&��4�tU�Tl#�PK   ���X},��j3  �7  /   images/98e5030c-de80-4894-a887-e6b61185dba6.pngջgTS]�/EDQA@�Ҥ�P$J��W!�Л��t�$t�ޤwBQj��H���^���ow����r_�
9��=����f��I����� �L��K�
"xJrx�-)�������#Dɂ��k0o��u��� ����*� ��|h��^���e�,���
�?J������
���(����O���� 
���_������צ�涎�v���[5 �������Ά筙�;sW��i��B�Ks�[FWk[G����= �5�1�cƿ]p��:�j��v��<|<|��o022>w0�B4^��K܉=�D �Cxy]\\x\�<v������|��@nG7[�[Wn[G�����掦����-#���;;'���������]a�5����ȋo������O�x���5�����K��=��`~���ǖ�#�����wJ��;�������Ќ�/��K���c#x����g�y��g��y�Sf�7*��@ !��/޸&�O]���~�M~�V�{�{$W�I"^_w��M�R��2�>���ʊ�D���M5�'_�xj^�ݸ��	D�D�r �B����j�X�:�%`z���2 u�2Ƶ�]1�/8!�>�<R��Gw0at�X��lD�yt|�J<���ʦ�����������I���U��'j�7�x�~S�f**�8,0C zyorY}=:r�WR���yr�~�M���F�|�ß��lw��a����*�f<ƍ���m��r�
Q�,,�@{�����y�I�y7���\��@�L�ǡ-@GBHf}r���SlXW����:���ҊP>�5�z��R��C;�kd�� �b(n<�*��>�_e�J|K0KjW��l�+l��%��j$�8�����=��e?#5�S�Í���a%���ǿ���M<���$�i~zr���!E���%��J=�R-�����������|�N)�<�E���7����gE�çtj�N[��қ�̪��&Y,���+��{XU"`��pM�E���]KB$ė3�})0YJ�w7/a�w@�j�W�󵋅e�=�JR��~7�m�3�P����m�S?��.�*ԓ-yZ��_i��X&��� I�>��IQQ��o�_�ƬOT��z_�u�ᡖ�܀XZ����_���5!���
���=?�'�I�V���?=X���ע������̲Ho��ZN0�}O�ι�@�D*�K����s����/$'$�4$}�Z�>�?_�ȷ꤈{}��Kn�V�,�I[���2��[�~�-�`�3�(�L��ć%o�p������7�q�2�md����Ϗ\��9�YY���w:��8��L����#+I�(J�b�mޡ��Z����{���
f_�"������B�2�N����k�=B�f �q���`:�n�'�3ht��B�v1ތ^��-�7UG/F���,�-)�ʭ�J���c�H㓻]V#��a1E�u�s�@�,9���fʅ���A2��A�.�Y���9�-b�L��x����.z�=������4 v8i:d�q�S]���H9n��$,�gc^�#�v���[S"�Z����O�Ȗ��3�y��L<n�6�j����=p^� e��*�V#'r}�G��ư�֠�9�\4�W��#%�I�H�x �&3���9�����}X�7&��J��{��G5�'Rl��j�y�����cy�m$�ªZ0g�����>n���d���?p��쓫�MCʖ����q����=��n"d�Ȩլ�R��n�����e� N9�+(��0��9�Aţ�R���g��k��'��A�F
������5p9���`�<�eD�N�h��7���̆-�@�[���h�r�]�B��ǯO�`�\��P�g�P�C�rLZCR�9���_�w����7�B�ڔ�+~�A��*�Z0|��*tX�	�� �� ��~�V~�b(�Ӂ����Ӎ�=�-&��=��ê�hy���9��?l2�� W4��e��4�J5x*�V�n;ˡu`ҷ�Iuɠ�#wK�3�)߱r���L�:��5j��Cg�*P6�>i.d
���	�k�l�B;�2ⱌ���,�߆��P�i�l��X߱Xn}��0����4i��
���Cz^�B�<�+��*��K�J�{�u��;�����.z�ڌ%���@�Z�L0�n�N�J�e �_C�L=�c�:�+P5��o��=�T��~�=�x�$2����SQ��n�6[���bms�/<�؁��o޿YA=F� ��5����C�VGBY8W�<Ȩ��MG��{���{���9GTL!�l͜�0��4� �� ���i�EBy{L���Gé��b���Ji�j�Q@!/���|eᙴB��� ��$(+gX��ܘJX��Z�w�ҁ��g=JZ�H�5��X���7 ��m@YGo���ٴ��2�̣�CL������&''G
<�/C!��w0*)�6��R����)�A�	n����?�h��������gFU�����`0w�A�$���t�u��&0UV N	��$���/���oc�G־&�5��%7	�� �/����t����#�rss1�s:��̬�����Z-�xB��<�|����RNC^Qq�d|y���$cocJ�҆s�?��f_" .�w+[p�VN��AL':e*M�cM��u�sβ�>��a�IR��+��	��ɏ#�~z�s�+��F3�\a-+��@��o/K���z}O�8���.t��u�p�=|�h:��Roϰ�`�����
K1�����L vL ��ɵ�`�N������7�����e��/넂��4����������L ��MІMyN�:��u�AlDM�><�����}8Vm���">��M�����lY��f��p�-�����F7��z�]웯�E5��V��#g+r���߾ڌ����O��xLr2�/B-ڀj��h��+�l�K}.{CY6�c�����l����Ӹ���{1=\8��w)��*�X���	��~�;j�$A�.Y	)�sn9%����������k}�"L��U� �+�T�2�i�[��aP����������3>��������c���=#�*[�yT�'4`0ʼ�4�u$i�or���Q`m:P���T�?c�����o}�q��̂[�2���S�8.����g���oewV�d1� �(�����!�m��X'sh�P4�q��\y�}�e��G@ �BjQ�H�$jӠ�HNjd�&�\�{��v���� ļ�.��p��tYڛ�J#�02�qsE��,�&H*�;v�B{�%��H��>�u�l�{Y,d;�7Q�I־?}B�X~�������4�;K$g�A��:4N孞��&���0�x�ؕ��	��!���s��=��+*g���\a�� 1w����K�4%hr�+3���ݾ-���1���j�W��ǵ�dw��Fb/ޒ��?�x�
Pr�lB)5������I��{:!��n�0s6~�q�m�b�}^b�G�	~��(#9E�t�w��ª 	�ׯ	�&���.�P�&˛]�	d�:ԛ���l�L�#D����g[�����l�s���Q�l�[M׽�E���S�g$��LT��d`��>w_����P���>�m�2�+�p,8s���-
��y\�t���y�se�?~�����s��߄;��R��p�'�e �Jh���}�7Of6���@�)�zog����͈�a��G�x�Z��w�õȠ��/�i����f?�SD�V��F�|8����g��Ф���ݰ��n�E����.Rk����8;�{_�CzA��#������r�:#�Z��&�����Ҥ����sT�P�k����]ѩD`�N���Ox<�ReR	 R���:��e-�Q���c<����44"�����Z�〠����޲��ho�f��ۣ�]C�~_/1m�f��.�<�1�#�'�t/�kO����!��� 9w&�:�>-z��%	�8s l���ŷ��n�������|4T�z�Œ��`"��sm���J�Ѹ�̱W��$���O��^�͛h �`Z:HT��O��RN�����v�rR�P��2�R.����Aw� ^H�'"�L�Ʌ�� ���͢``�ixTS�;t��|�B����<���{$�4x�V���(�����T
ŋ8ѐ�J|�u�
	K�������:���@��ʞ�3���V�]Tr���|�¸9�%G�k �O�>���v�X��m�v|�qx�U(@����x���D�(�-X
�7�`�`<?���,HC.yLd�c ��D�8,z�� Rx���G��d������vu �����}��9�'3(N��V{EY��ss��9��f�`]p��kӮ�`O�)�t؏�w�u�9�YSu>�up(^{^�.Pdyv0�f��ҿ�,v.��v���T8�f�M,����'�8�Ӹ�/V���N�j�����������K�)0w���t�Ϧ�������(���f�y��W�6G�s�~��c}ĔG֓����Q��3��:��q:������v6�H~�d\����r�ז����m�D�D�_��	�}�/{�f���B46Z8>�����|-�ц���D���tf��NF�63�9S�}�W}�6�4��i��~�zၼL-&��9Fx�gf�pW(� �(�L�V��7���7s5j�rN��s;�f�+6�6�><�(z1� ���\`4\�i`�r������᳋�S�|��H"c%>_Z�m�����a�Z3	�~Byd3�w�U�W��j�xD�eN}�U���3�SudgGF�QČ0=O���ׇ��Z".D��~m��N�قksS1�3<�MәM�8<�c�,��k<�"A$v�e�����y�a�p���d�1\�óz�	��X.�ļ7�;]WCx��ǾzjE?�����������=..�V8'K��~����x"��W��2)�ƢAn�P'1	���U���tN��H�����N�k�*�[�?j��X4�SRt�op/y���6�HT��YEm�f��Tj�w�&*O@Ȼ�$<m
�9�7/K>]_i�mbq�^�|W�
k�E�h3��T�$�Dke ��0�d��4P��{w��3W���s�:"&����h|�W��_�̶N���0��d�o�w(T�6pW������Y�.C�H+Dd��z��_�d�Ӡ>�.�b��Y�k�dP�����cE�e�Xc���5�/��-�o��<b(5�[yֹ�g�#Cξ'�H$���\���7Q�ǅp��f��@�������5�&[_�����K���}���z�x�����Ѭ�b���a�\Q_��ۦ�A��Dʸ+.$"!8���{m�=PsM4ԍ����Q�v����TwZ�����998Q�? �&g$IZva0�{�W�l�l�:����Ċ�V�P�)YD.<%���~��N\�T��-h���y��Q�Kt�����
�|�ۭ�U2[��� 7���ö{	~4:�����/p����/w���*�L��"G*����K>R_����1ζ5��+�E���K����뽯�a�y#3/����H��@�.o��6q��)"�HB�q�lp��ѦvH�5�d���Ö4��w�I�~�+(I=�輗1�I�X�N�?����X%6l��?i�S� ��gʸ�{�t�V��Z\-�ax6���P����QnJX77G�a��ū��}���77�����	��R0n�O^�w�_�l�c>z�ؔ2`Z��&�0��K=�݆��4A�����.q73�1���	�}+�o)�B#15+:�oM{��{���S��+�e)�N|؊�v�8�Y!�����{�7�a�M�g�c�۵rׁ=?�	��G�3�qTW���-�"!r(��E���iY���'ι}s*Y1oLT�YI�'~��5I���~���+a�X1��q�=!1�T	�:n���,�����+<�2}ٿ�<��XZ���=k��8���2��R��N.�Tk�uW�̼,y�}\Q�#�;�'G;AU'W��*��XU��[e�Avٸ�z�)[�U<L�<K�	�
���A��0Wxz���u|.�;L�L3	8bg<�b��8��+�ʟ�H�H��̟��F\%����+��_�_�ӆ�/��Z��
�6�j���_�?�w�K���;��Hl��$�=�z�K���<\�״<�d���a������D�f�e@�[5�̱��IK �骐�?$'��6C��~�W��[ze��$=�M�3�s���X�f����|C#[7�q(��!ҿN���ԅ�~���1�p�����%���ᝲ��+��[9��L���Q`Xi��؎���ϥ�k}_���d�g++"ifO��=���5����y�����A-,��L� �í�{����f��V�����ƸU=���C��QC�Љ��>1��~@�,���F�ſ����sXX1����9�g��D*��� �d}��Q�8����?>�H��?�����1�(T�-��lN$l�+¿�6��_U
�;w���ãӔܬ��@|��> `x��a��
��m���sc_9e"��s��.�V�]�ߺ~�T+xw�\8|�pQ��[�w�����Ӄ�;y�^�G��%�{�z��p�b7ٖN�5v�h�������`9.C6��.6�9��ŪV�~���`y��3���ȇ-)>������'-6vnb�������X%)�����o��&ӫv`H�QK=}���C�4t������9ל��ӭlĤ[�(<V�r/}�7C�^�QF+K&b{du/�iA�<<2LAng!��l�I�0>�����.����ݨ�q(�/h�u4Vޔ��9Z�K�a��Y���~��3���a�󊕖=�~\�H�Q���Cg�6�,���fc�;�n�56��^��ݕ��K�sƐ;�\O3���nn&|�WZ���	�8���p�U�����y��S��K�3�[��M$�U�7厓�Bv]�5�H���M_�����({��P5s�a�0f%��;+x�6c�E�l�Rivb;���N`��������+t_�Y�]ݠ�����80X:�/���C?�W��?)�֫�ga~E�q�̠����S]'�X�6��@(؛`J�,���R�:��*ݠm}��7��ӏ��G}"���'h��S2#�}d������z�@r$}D�F$`0*�A�)
ki�ñ�	�)g�ʨ��v�z��=���=Vn�+�a�G�e�|}7�m#r�q�W�r�H���]4�X;��^�*d�Ut.�he��Zvɟ4��ڸ:eS�٘�hU��}��[*��5�ul�i�wg�٧�P�Z����kY�"YE���Yg�ΐ�j�+�sm_pK�F���<������o
�T�4H��:.�X�C���*�Z�/��qqN��:��Ĩ~cH�6�ѣGc0DO��@�!;�_o����L��!�9�vDچ�-k��8*�|�91�I��Ɯ}��n��&��3�Ξ=H�&�bde�cSe=�#��^��ݮX��Ǫ��?�eRc�h��9R�{����{�ȠN����0���6pX!=%hƨ��=*�S�׶�P���K���m%����e���nq&i�~��d�}ȡ]ZھtEl�r!A�\-]w�v� Z{��QC}~�U���h)��;�7!!Xbʰ�%yZU��R���RxpT�X�D��!������(f�Ѽr�����Ə��Ѹ	��Ɯ�>C]Z�DRմ�8���A��]vc����8�;1K��jn�e�Qː����:�2��jƖ��	K+Y-�"Gҧ����O�*{H��� 1	�[�6w{��%$�YAK ��YUwύ)'�Hi\�Y�3���<����ܧB
� ��5�)ٰ�u�Z�>�ݳ(�rP�Kߚ�ӈq�w9�<�^��E[gg�υ[�S'�#D�ް/��ĭ�����I�ޖj��8���ʷ�g���͂�66�4pk�]�Q'��G?la<S�)�S/99U/S��.�������Е��K��gr�xq|�=p������\
s�`PC�kZZҰ���dJ����p�7vs%�c��D���C'��xq��G;�ـt\O���.�V��~�)X���"ߤPe�����r�)�N��y2�/���u��
��aU	A��L3T��	F�ܽ��iܰ���c�E%�)���6�<���~��>�=����[5�c�6�8J.wn�?����6�8�Qo/(p\55ɓ@��W���I�
U*藻���dD�ߟa�5<�s���+X�t1;,�J)Ӱ�34�'�>���fnV�!�'�4Q��p�:+��:�ld�Τ�R�W8�L�	���������T�b��8����K%����U_c��\�%�Lom<�n��)�������zϫ�$�o��k���~�����RYͼ
2Y����MF�f����6X��E�Wm����c׬O��������c{�)�P7o�@�=#��p{Q����?X-+W\�� zD� ����*�?㮮��I �~�{O�D��ё��">��e/Z>�,kSQ�FWZ�<	�D3��.$���5ƅu\���>����P?����#pl�������M!�=\���P�Z�^���>f�5�)��ϝ�Ie���A$�|�2�Vq�ct�"�F�R֔={5@�Dw�+�5t�l8���v���k�g������i�T�ޣ�'j����d'4?��n��k<���O�c��Q�e�~I^Ѯ�ث{W0��Vm�f�;��Ii6|���χW�w�p���.�<.Ɵ�8fX2�zkT�THW2�;�3r�;�~��[I,.�MV8�B�̌v%)�^y��$�5�r=�xq�*�?���i���}���<�Q�����/�ٓC!A���]ݜ$���>�a������`�G��& �;n�x��s���e!�����������	-H��� ��Q�3i���|�QrV��MX�Rq�b���PN��%�rS�G��]"]���m���5�{�d��9p���;��3 �q�����IQA����6��;��t��YB+��Ʃ��b�O�0rCG��1�J�ƍ��=�mĪ� �ӫ�!>5�ㅼ{��/��הN_���%�^>	N�ak�/���1)�9���63�����;����P�q'�<͸�!�߿�7asdŉ�@�M��s�*���G��S��(��a�
��jAh.��$M!�~F��c.�B���=�A�)I+�K�mš�Aʞa�ge�pW0.f\о��W��З��s}��5<?�K"��4�|�[$-|��]n��zC/���<"P�!�i����� ���D�/¢�+]�N��~)�șnr�������]�Kh*�G���oe� f66E+��DQǶ�Zyo�#>}"�yk�\`���zgT|�@;_�0r�̢{0S����g����i�����,�� ��onj~Ybs��缀���ײL	"v��aתr_gӄ��L-���9m�"�LT���ҍ2d�j��28- Ɨ`���E�8.-�@h����5��G^����g�����x ���M6�'U>�3�{���/��RM���6���D+]Sk�����z����se�������2��������y��V����s)���VP�{澗S���9;����t�q1���d�\�����b%��>�!3Ǘ찿����+g,�6$Bb��/�4�y� y��2<��s�ĖT9�S�v;LV��4]%�w�#��:��/��DζЮ�*m�V:�,܌�/��w�b	�j�v���x� _ĎU/�C�b�iz�*���ŏR��6��z�E�,�)�]-�,dy6��}ۦ�+k4�A�Z��m}��_z�S���O���W��2�Nlg�D-L)�3B�'��޺��u����g���Gűw�U��do �	j�2�"���{�̙��K�Z�E]}�%���2���w[7l��aAa��<x����b�^&�������G�v�ĥ�V��zN(���Y�n$=�KƒH �e@-+e�``^٦��WȵwS$��ܭt":��8��La�C��N���Ģ@���*�����y�c̛����7���.9���6"�$�]���(^n����&���ܐ5K���F�S|���czL��U�qa�䅰S/�	
l��$b)``utؠ��:[������a(�ǣx��:�����.��]t�4���	jo�r����(uF[_������)B���WlR.��塱�J�=Q��g�.�r�X�6����d�oJK̄�<��v ��d���qj�o&���\�1���RQ��Pb _�c Mno��"e>^!����a�>�Ų��l�=0���G�=�w� �1������mGdC�#�Z�>q�J�i���$��*�a�#ġ�A�����%��^[ȍ�!-y6{?��؜sV�7̱fV'S!��ki|Z�1�̸�x�A�^n���i4��F�S�o�����o04�]Y�nɓ�V򩕸����(<h~ϥ`Q8�53�F�?Qi�i?�Vj�KF� >��<�u��T��=TJ�'��b�����#\9�8���=�����͎wj�IRWG����D���!>��Q
}�ng�1Y#�p���`}���Ӌb#�̓���VYU��^#�0��J�f�l�`��Ţؿiya��g��>�N����k���<A�{Ֆ�G{�E�F�&��K2�S_��gg�z
h�o�8HL�/V�����	�1�^�*�U�Dj��q�����>��-�?ɗ�����ЭH!R�O[���g�W�(i$>����@DY�~U�����G���Fm�lc�?ɼLx�"i��,�,+l7�6�� BAŃ�A5��p���ǁ�n-"����KOO�~m�lU}��de� N�+':����J���Q���@)��e�~�:��r6�wB��'7����&�D+U����l�<������E�GË|ug[>/�,t�&����+���5
�kݽ$П�TU���K�xсR��7zLƨ��A��=�CUq��oќ�����H(+����!�L?�]��|y� ���� �Q^�x99}Ș�+��?��b84����f��G� ��S�%����ӳ>3��n_ڹ�ku�1��STR*G씘�3��|&���ӯM�i�1H��*��1$Puuu�B=!E��B��z�%Yy���U��Z�� �ET�����6�e�8'e���3g�x!�i�匇�����j8
:�@���\��p�Cr(����;6S�v��ݶ���.3�ٙ�Z�=���&�TTl��ة:�%�4�2���5��-}��Q3����n038�$K��K�N�#j(c��M�5���ksn%�LGlϵ�Ѽ{d�`���|���|E��گ�9"6��'}b������N��JN�5c�\�gs�v��9�)">�_�`�Ǳ~ @����_�:����DU<�'�^%����' ;�o-d���������>-\�4!"�,�e�mV�f��Mb�������D@���p���ށ*b%�pyq:�!G����CF���?�}��x4d!Ƈ�G�+�hC�Km�,����{���U�a�������tu b�������!��A)��.~؏�|��w4?��&bu0�ڕ`��A_g)E����~=���Cs��V�8s'���%�Sm�j!0m��/G�L�8��������&2����%?;0�z��Qܬ�b�x��-��[�òȰ.���&������!E��@��K�f_���_�r�Cq��߈J��L�bBP�o`�e�D�ϪO����Igk^L�ꬷ>dX�L�#*�����Z����؎�^�8����ꧦw?PʔY���^u�]�/��G�ѓ7M	�l��JI;}��D�񐨡\/��	pc��C���+(�,��/�{r^�)&Y�20Y���ؾ!@�{3��!��2��e����Έ�ݱ�j�/r0��[��kk �)"�U���c.Td��Z��>�o�m��U�R�F?���Pf�+l3�q�����/үRi�S�6������\��8�zK�+��{��,�dш�r�Rr�Q�*��N���|����R�=�P%&��Vϐ�<�Do�ݸ�W: 2�pV����D�H���u|Q�����3�̔4RPU��[G~q�ʡ�`4��j�Ȱh&|�Y�icr�	�D��KJ�PY��^[8������`��Y,|������[����υ�i�m����ƈ�|m������_eHG��b�U������6�d�Ar@�&ڃb����#��&��{��5��
�������4�=r�������77�6��  )ɵ!�fGl���g]�����I�=��_�V-Z�xA�ne��A��������ӿ�����jX@#��c0+5""B�۫;�aT��`0JL���\TT��RC,������
����o���J	����Y��
����>_@-B� �����ڧ�?/����z�1�ԝv�u�6���i��d�wLxo( �ΰ�1�Q���}�٪)���x�,%j�ㅸs����T�2.i���B�`�FKky �I��c�gW��)�L��]:� �m!���� ��4z 6W%	����:T!�Y	�7.�I&�������[~��i����ݑ��\����y;�aX3�\Yj�~�m�N�#1��'��އuϓJ���}u)��<��i�p�P/S
F�O7���Ms^�-޴�����Yg6��u>�� �y���>Z��D+l�8~Lnj�������;�,�:�3>��ƛg�ߞ��%)w��냵1&�[�2Ʌ���C�/hw�7�~�lY���/L���~&����3Xp6�ȧ�7�TXi֬WN0��٢ϝsuJ�?]��?�3E����;y��ER&��PK   ���Xǐ]zd� K� /   images/99ae2b82-1d43-4592-a023-63b23200c4a8.png<zUT\���n����6xp'�C� �� 	'��4hpw�����ǽ���sN��N����]�j�WW���I�	  p�e4  �������u��Bp��$���< h
2��^&'�h�����*kE�g3"��n2'�5�k���}��z��k��Qr*��zQ�E���P�AU.%}�����	�;ޓ�k�EA�������5��Y����� w�+H�UhQ`�����	�dC��_'$�Hn���o�)B�х���Զ!b�`�[�������߰5��:�r�v��khL �t/�����v��K_-)��i7�8yol&�ө�������;�FF;����d�^#��D�a��|�����i�2���O,i�B�K)����SJ���	�d�`�-ǺU.��I���_�a+^��G�+�X�Ǹ��K/R>2��W8G��R�%�.��*ou�G��/�H�9u��{<i��'�G���'�*KR���k��n3V �6\�;l̊�n��K��x9���r���9�/�J�h�~В,y�t��J����L��H"ˊ��r�k\�}ff�ƟgVH�a�
�q�,T�l_V]z��)���<�#=�B�6f�z!�]&�5��.;ޤ��V�������r�{�n���������)Y�km��~��$�� �gz�����̸YN�#�f��x��~z:ٞs�t4hӨC|rS�ǅ�9?�UFr��?M�?����|�>\�5En�$GF]��O�=�_-;���>|֧=�!�����X�38x߹�s����SǮlћ���ۂW"K��� �r)��pﺐ�9��_��vw���ֶ�NW�Η��G�ZVe��?����Qۅu��|E�켙Qz����̮�+N{�%��U�ݪ͚D��L���Z"k��Ǆ�J��%�k���< �z1�*���Jy��DͶ|Z��1��3��
�ٴ�d7��[�7�s��y�j�sL�kH�\�o���H8��t:�5<�+#��6?̮>`�H��&)ο�P111�WwN��ڧ���*$0&}h���:%��d��d��۱�5���a쳨*����'�A!�+��G3�)�t��]E�0G�4|�@�����]�=�'n
3ާ�����0c�oi�-3g_����Y��8;q�t������Bt1pVc9#⣙�tӷu��p&��������(w6>�T��i�
��i�|4��@k�lHش?m�J���敒9DX�\N�(�
<B��T0�+k�.e���3��	��!���*���l������Fυ���w�o�Yz�]O���)3��P� �������Y�E��a�k���VUq��in(��L1q=�5��s��,'{1��L~ ��d���<m�t��n#���y5��ξȸe�N<�B�x�h���0M�}��]�C����4�|�ʯ�;~�\���<"1F��0���(����cCgK���;cqC�d�����5IZ�ln���_�Q�����Wnr����Y"�ٞ=�%���������g�)~-�����O���%ȈA�����cRdR�}t � bn�����8U����d��>��i�����IN�_?!�}Â)�ӃfN�j��z��{	�E/�vj�-��gBrh���F��FX��AꜾ��h���G��I[�l�Dds��if+�Ṳ�q��>�l^kE/ݧe��>��߀e����·\\�������<�!���GPeG']4��k����F����?TE-ݐ<8'k+s�0��Ш�����x]j��U`C����]�D������/��M�'��⚊�y��26\U���~@
ش�+K�S��CZ[w��`n\���p�A�u��h�x��fcƷ��_�c��N��!/���*~G���Le�Aċ��
2����!"�0m�Oq�ّ��o�v��'���=�r�1Fحt�i��BC���يO��]sB����n��@����1��VМ��K(�}������	�}�(��V���%t�p��UI'�^�P�7-��K}�:>bk������Z�S�W��T��sW9}���}#�>�~�����Q�bР���bBt�rF��Z%~2�c�����������B�!
ؙ��μ��pu�S��Ɏ�PF��Yۅ=�5�[�e�J�$����sC�(�"�tc��2'v����%�A$d�9�z�����w�TmE��꽍#�)LP-��>#��W�.vw6=D���
	~ �l��"�n=w����p���Q��Q,��j��LK�7�vU�6ϔKX����{�����3fݥ�VH�����W�+�s�ȵ_G���fz�+L7�e�8�n.�Ґ5�2���#Λ�N&-�Y�P8�CC�g��|-:_,��{���4�zb�Ð���Qң��P���I xP��� �@��pR�=�� �Pm�3��|��l�Qd��5чV���A0�}�v�{wS�� ��jX �)�s�e��"E�"�����kF��/Oi{ �n�*$�<氿>�O��4Hg_!1�fc�U�8�c��ke�R�9)y�(�6N��T0�tUi�ܜv��]�e5씪�ٓ�f��%��,�b���Ǝ��/CJ����zd�(���!=����*$�G�kq߄;����s�r� �QZ�V��]��zE-s9��8���ɛi��侮��չ'~�A�s3�TU�����#�(�G)�-�K�=�m	�S��S5u����U�ܮ��T�}[n{���H-�Yc���~�ը��{�����=����\�����3B-����RNB��_i�J���8v;*k��g�ܶ[����AU;F�$]���2��.dA`�� s�w��8h���~��x�~?Z@�뚸��\.�pD��O�����h`���@��X�~J��K����|O�_�᩻&i�1d��>[�7�:�1�6]�bW�RC�E|6"4|���l�tn�#]��u��J���o������a5��/����o�{���-i�{nu]W�; �z<	���_��(�֫���F��nM��d0��۵�@ ����ˁ�2�v�t�Oܦ|k)>��+4� ��=��o�/�%��~���[�92��/]/{N�ק��}���ވ�&���jwP
��dm(�AN���z8����%�Q�Aܕ�����@�/�U�s��D���gK��N�����WL�G��un���!���O�U��f6�2�*�?`�
ui����^�q�*_���ٷ� n1M�	O�����Y�|^[��~�R���_1�~��~��|�;��bP���"�g��訬��b3,{tt��� �O^)1aw���rнvZ�q� Jʗ�)�5�+0�n��y�4$�5���Ga`�Y���H
e�5F����~<��Z����s[�a?����̴�P�^{���>�r4�]��f�+�l��1�tߖ��o�W�{q�����0�Eد�?�$E����.��;w5�R,8'T	�?qepF��zf�!�UX.�i]Ͷ��S�/N��{i�����Ǎ�����sEc�7Za	����B�	O͐�Ւ����=<J����fE���s*�U���2�
�'�N0���ߝ���m���A��՝~���~���ߢ~M��ņi��j��LŊ�k��x���f��{�s|s��Κ&�K�-z�$/�g~���T�5~*�+�gr	����>a�܉b�*��M�J=�Ӊ~��^�7)z�f_��$�����5������o)�Fp�MQ��N�B���u/<��ڬ:z���='��?���J&�:��8����U%���� Oc1c]�O�z�h�/��LŶ7�h�\!�~�7)�II����"�����S����y�J�M�`���]�m�MN{�xh���Z�s��ƚ�u�������/�D�r��s�2�`S�s�7c�>�	ճ�'�}S����Ӥ$�����J���WLV�����5��t�����K���x����q�kd8U��4�?��?�O��¦�T��_�L�:�,W�^��l��H`T�3��P7d���3�����(��"����N(^��S�Q���+�K��������⼋�Ѓ%��	�y�9����݉���~�}oܴ�&k�;\$rw�J�`S�����A�ۯ'�u��n�|^ú巏�㧳n�k`�'��S6fV�x�M��� �����v0�ړ���*"�9��
ٸ_��`n���9x~ �e������\o��:���7�%&^���k�?�,܉V/�B~���Ia�3�q�=N ��t���=������-�dU�w�$c%���>~���O����c�)�#�O��4���w^�H�R��I�Jq7�@a�E*o��u"�E�F�L����̬m���M~���;��J���S0HiJ�2���lB���b�����OW�Lfz�g��T�m��ԏ��	������-����;��Ґ�(H�I`�.[�%���(�<Pr��8F�"01��>�/T�PCS�:�b���(x��[?��I�������_��5O�)����� �=�m7��H�y���c!#�Xm�p�P7<`��EPD�����Cm�?!���[1�.��^���l����p�6� px:v�ⱡ'8T�,���r	��X?b�@��@��&:�̛�L�*�׹��4�J�e$=�{�
:~|g����|�!������:N��$a+�9������*Z����j[
Kg�����}Eze�j�lM������B�Ϝ*�I�@=��6�/�N���D�W5m�}0�� {a���W�q=?eHP`9�!�����VQ�?����*rJ9�q`O,��L�H�����������K�ݱER�a��@r�ȴy��P^H��`P_��u�������I�U��bD@?.��^�Mv�wN��n�p���[��a,� ���B]X5���?�qzP����I���m�wcK�lE��5���OYh�,e:+���靏b�HA�^eo���ybW5X�9��YBޑ��T�Sb��{ni��z�p_
R�o�4pc����i�Z,����`v�d
ėbv�W�!�4�wj�N�*���y���3�A���[�/��&���fX�d�oC4�
���+2Z�B��$R���
 YSu��P��G��L�m�*�+���mVp�]V�ix��%`�/�]E�-"�w��M��< V�7�ȣYL��k0�P�g#��ڌ������`~o4�c�0q#Y.�4z�������e��� $4����㪙��f��zǕF�S6E�)�+T"?�Sq�P�ߚ�(��l�j�����{��w_W  ����K�ru���-!fjm��18��="K����ڿ���Q������k�uFDgD���?j�KmTk$J��	α �X�����$5�1,7��~�����d��]k�����)p�\�n��.������F�{�jƎF�d̴���mX�dvg8�����3WHC__!�ԫ�[��[�	B+>E�2��@��3h��5���'��f�}J���zF���6>/M�9�ϝ��^M��b����[�j9��9-��*����Uʥ�+M�J�m�l�U���&��7�䢺����P�b&�.��_�1�N�y�>\�z�9.[	���ǫ�K�<�����Im��:�m��?�+#'?Q���ǟ� �J��OXgv�>���{9��=/q%l��C�f�:n9�*)&]��'�j�LNz!Xkd�&me�<Ԉa�J���O'��O@��4h�wL���ZYխ��xQ�C3�.#QT��R���ٚ\3	\Ԥ���ے(�����_�h�
��}c���U��]�_���Zj~�jr2eec+��d�B�:B���I��^�$I�#� �N��0�fe�q��gOT�U6���� �f��]ۑ���}\���b����:o��ɗ���fb���\�茆�ژ!��Y�x�������P��?8����nch�i"���շP�Άh�'eP{��̻����{8i�wa^�b�qw�vt gls~n�����@�7�JƸգH�_!�����t3�V��Ȏ��T���|������� $ ��r!�8����Y�X��;�7�2W"*���+]�Ի���2������o�P%����C���ҍO���6v��V�)�	����X�$��w�<�l�/�}��h2ǟ����ӛ}�K���	��Ҷ���]�(Wgf������Ѓ�	�zmmu�%T(����F�sY1n�O�+hb$�$Yon�w\2��Y0��r�9������=m��������h$���Ğ+}���ǭk�z�Y��Y�+Ĺ&5P:���H`�%r�|��%�sݛ�t�gw�i㊗��]S�t�B�A�g^M@�'��@T^$�_�l� �x8=�"=M���w�%Z�2�Y/��O۩�'u�:V�2�U8֊���c�v��C[Y���:����0�����Xшo_�������Q��<���Lhܦ$ad�{&���w��E�<��*�!H�u�|�^��M%AH��7gk�8��%{�� �o�̸�)�����	��O�	���	����)���@�����A��A��kD��>�t�m �D��8�A*�m&e�J���<��c��U�I�p'<��]�+�Y.ܤp+����MB��~���=�cN�3�������m\�lkB����W]�ǩ�P`ӼC�gЈVֽ�&���b��p��.�<ߟa�/ۣ�6a� q�L�o�A�L�^t��y~��e���������?B���:��?#;
_NS4{��/)N׫��Sl�f�'M�2�X����<!���ݻ�{�F�W���n�'6՟�����6�̤N��t1h����e�j���^�d�"r`xC=By��K��L|?s�����卟�h�xPuR��r�}��nc�0;Y�m�	!8�A����&���O�ߜ�)x��!2�:������=���7{P-h����bШ�h@41+��	`���}4WF�I��k�!WhS�L���}�9��"v�[��m���Q�6IU�m�gY\CT���ǥ�ĬG�)B�Gs-�D%���єj7������/>a��/�:��uA��
��Y�3`%��Rc_�x�3{��d�Щ�r��p�i�XV,�L�ڨ.�[�n�r0TS���$�'�x�����]�	O��w�\v!�FFDx�^�͂l���|X&N��3���P��^|��؅��:ϑ�\ ������ �Yq���-����q��C�J�z�@�7�+&mk<�e0��~��t!�b.�OY����R�[̘z��p�&}RUm/��ҿh���ߟ��/I��_p3$��#��Z��&'p���ɴz��o�s"�X2�)q��z"O�)�.GP��X)m_+����'G�u*Tŝ�kHҭ��.�mȶ�nX
�gg�P|���,�%:i�.�"����i ���3��qS�W����4�R� �v���esCd�~��w�.��u"�=s��bv�NC�  �s�0e��h��˙g�h�� ���8x*���Ծ	���R׊�5��᭦�{1g�jֿ����_�{�Ǥ'lRc�z�#0-���Q�4�41~��-���)��.��������jFZ}RJuq�L�*`G����Ҫ�Վ���r�J���9�ի�h�������m)b�/u��.�<��6��2�BM��-������s�O���U���~��͙/�dyd-����[�Kq�mXM{Z�/�] 52�"�T��-f�\����J�k�V�k���U ��C88/u�H�Ġ�@��y��n�/��(�Hq�"���ȗY��ea1B�4lOeu�g�kJ����s��͡�8��"�5D�{�����+05�L>M@��Dy�e�l�I
�ȶzw�����A�����a��{o	�=@U'���Sd�^�����ytz_�_����u>̷Iw��mћ��܅
�l9O�sF�����|5�:���	{V豝�A9Z]Pg�{��~�C�Ƴ*������1����3!��(>��S<WcQ+q��c�վ.Cy�qP4.�x��ǈeh^qU��w��Ƀ�a�rN�d\�%�3�D��]��	� �4��fv��E�c��6�^1E��v�	��_�
�@���r��l~��h��{�Ag RP�~'�r��p���1*�W-�/
�(<Ȅ�ʐ~�Bu�켓� ��hx'S��A��6;F�q6�E��>տ�fUZd?z� ���H�E�9,�GE��S��$]/�Wd]z�{��¹��Ju�1�|�9>���U#��E�����?��R!v��%�
ٜ
�hE�"n�漱����5T�-�ٖم�ݮ,)J�ܨ:n��$�A����h������vK��z�GS��+&�J)������z�H�T-�Dج�4��3�LN9�u��`�y�
�>^P<�I&7��/��%:��F#���oɒ#N氎��d�۹Zs>o&�4�#�'A���)�f�*���#<�Ͷ�m�w����?d[���8��ƻ�U�ET��L6�J�D�:go����&��[����(�� �D�E����7�y�P��;�Ks��kn�m�*��r[Q�Q�"dH� ՙ��t�_2*(�:��z�n���B�Qi�N-�;B}�ژ� l0ZVnD)���
ǐ�2����[�;[�E�E�,D�Õr��,�%ܸUx%��&�H��:�e굉������'#�X<�7B2�����R����K�Xoo��&,�T�1(s�<�hM������+W!R�g.:�O���";#o�~ˎ���a<\�{�iP��ś��<3;�:�=��nzg8l�aC8%Z�*�ŠÂ���o�����4�&�·��X�*�㢶B����츉�˧��lo�a:�3 ����T�;�)w��C������R������y���Wg����.�n�&<�u�^���rr���zȕk�8�|S���/�� <�w�L�Y�;ӛZL�)D���k�V�����\������]�I��ӹ0a�t(��\�j!̾��\�x�?�G�i1d�T+(K�<I�,�i��w}���k&G&���P%�D�Z	��5˘�����g4c�<�۔c�;0)S&�K�;�����<���Q��ϻ��ZTt�]j��J���l�}|��\��UC�y�Z[�Kժ!�E�Xhucw4%\2#"Al|��ƀժ�.{���q�L�/E.TC�oI�Z�x�b:UQ�1�!�)�5����DšR�*��_�z��$[�)���M��1n������cbP��4��
h�����V��"ǜ�?}Ǜ���߷ߨb���Ԇ)#���j/�����ٹ.��>�����t����Ƌ���M��V$k։�$[8�#�7YYX�z��q�n��L��Ɵ��.�?��>B���s�8l\ϧX���ZBb�$�]�8T�nLm��'|~?�ʝ�K�����-��������u[�X�6�Y����[��K�m�$)��Ȧ[�'��c��cɬ8f�7A�W^�|��p����?"�WՈ[I�$�2�w3s��a.Xl�u���CPl鍍�[���͂Lf�����Px�Z�������;�4<q(m�o����+��%�w����:T��=�9J�4�[v���@M���Z�<+��#	�Y�\gzj���;��%W�7���v���Z�����gaG
&��o������uo��\�*�Ci�Sd�齅�X�K�x]~�k[Ä�������pa8��'���;����J]`�}pF�$k�aӿ�]�b&j��ZHJ����[�Nj[��{u{����m�s���N�Y��&ݙ��qw���x�2�Ѭ)��W���g1`KzI�-nzX���_N���-�#�?7j`��r�/[�D���\>�u��L�Z�13�o�B�9.���h�4�$i2Y���"�����,C�؉Υ�-"� ����u��p���ꢁ���g@�������۱�`�=I;���&j"����NmJ��am٢�2WP�&gr��#�2�D<j H�(W���B=]��?���Nf����/N;t�"���t�}�tOF`��S�+jRԸ���d��G�����i�H$= %Z�}u{c	M�0];RJzD�<S���u�v�Q~)gʎ`B$��Hf!��+Ֆ^���̠���_=��8ABL���Bq��zb���R�W�rImK��� �WpK �=��c��I$��3��	�Q��_���z5ʥ�4辉@�:,J��'&bY�A`�xr�s��sm�hD�&�+9�O����tk����q����Wr��`~��� X`������֛KS��������������)��ő�x/eV�C+,v� ���*S��yW��<~ �4� ?�$�i�C���V��w��`�����Ub�`������Y�%��}	H6��P����B,"�G6��xW�C����'x�H�T�����e��W�<7T�GN�����'[�caE~Ks�3�JGN��t9���3M�_Ռ�-�y�;o�S�������zC�c"k�%���6� �b�e��x\#�� �q�|��9�s�]��eM�fV�E�/��ą?&s��:U%0Q	e���F'�ڇ��U';�C:+��wބyMy����*Y��|ǫU{L�e�,�9e&�n��«4h�&�4Rݴ��&�K�N.�%�Z2����\،�z4G����lk/V�E��e�s;�
U�����du�`g�sҾ�$�9	\�������beJ�P;ߣ�aml�P�y[�#��������_�a� ��ƶ�s���� ���n�
��	���nҠYD�OY�aM����y���u���>��f<ݽ	N��Y�&�����eq���{���9O����(���&~M�� �Ѓ!��?����*��!Ѷ#��!Q����V�C,H6�7���0]���ϭh�h�c��9���{N����?�����h� �z:57Bb�Dy�D_%�8HB���Ys���ęS[JsY���@A��O�^&�9�+�k���e��(�n߹De!*���-�a��58��:�C�~��p�fiF�1�1�1Cn�������DJ�m!лTWN'�,����8�>���A�
1����c��񥧧��f2����e��I��������"���=��!�� H���=c����rj��,����|6m۰�8!\˱��Zo$�;G9����mmy�cm�^�QgHTxIƕ���N�8	����˭�Uܐ=�N�>le>�|�i�̀�ާtt�x�7�u�<�o�es���"C5>��h�c1"Vo�l|M*��q��wk`Q /-���$�y�w1�@�����Y+��]w/+�� ,��s�׺5)�}5~T�a��i�o��hH����?�b6;���OL��5�|C�i7X�<��Ϩ��<���+?7�kao�`D�)@Խ�ː��l�?׿��G��_֎�A�PAD��Hj�#-��-�xi��3 �'�H�H�Y�-�"b6�y9@��=��zW�A[O����P{f�)���*¯h����3�B٦_)�4/�E2m	?�M2�h�#d♍�L3�����G�7㏕2P~.�3N	E����������ܝ�B�y����yO�TA��z�/&���BP�d���u�;`v_7]|B�I�]8��Xn�2h�87�{݀�%�]#��;�����ʈ�0bA�� ����#i�a���D}?Gћ*ɻ>q4_j��^q!��?n8x;WR�@!o��(��B�Z��hh���_�|��§r�/Y�(\���i|���S#M��5��O#m�@} 
ܠ���E5�������'x��\���'�y��̅y�Ɠ�ѧ��d�>��*���&�Q��tI�_1���3�`;������B(�:Y�P��`�<[�NŘ#Ή(��op��Ѥ�y��M�M%�j�w�Xۘ7֬`����R,���/Uk��0z��?���wD�0�V�~i>�"���/W�S[�?V�DHBzs!��5�(v����\������fDh�PG �������xۙ�����
�WR�+�j ����x�Tt��p/�$���������ĉ��;	j���j �⎸���ƊweI����	��k�X�13�\��ݓ}�
�_w_�����=���HO��m�v-�S�-�U���8I�N�����Ln�
ɭ�s\d�ɸi��`;`�Y[�Gji��ґ5�*��o�!�C��)�������p��a�z�Jز^%ʔ� �� �.��;�X�I�Q`�G
�y*�xf�3B��C��@���%"�<>ܜ���7��MƮ��b]���o�m₌O�<�A�@�g�Z.�u1z�����D�΍�u�S�fo2-���I^�R��t��0��M����8����H��h�ff�8��<�M���"v��Tؠ���f�����z�՘C��Dٟ�xɡ�oe�����paRD��W��1m�����* �k��<�.� �wo��.+03�W���[���bUQ�g��,����T����џ��l�-�+P�	�x�Ar1ЀBc��1���ˏ�wJ�� p�oN9+:@���8��RKbBN7�N+ӿ�crrO��[�=.�w��d(/fj�lV��&X�;�ϱ��ຉ±��@�;�D3Y�bCY�L�)��@Pa��6*�S��[d=#�["���R74�����&�֦$I��1S�d��[7�;t�]t�^��7B ����q��u�N0,KS�\�X�(�8��C�q14�*!�B�^Ϧ�������ę^I�~\,ߦ�Sǀ |,l���[��!��z��[ɲ��JS2��Ԩ���L�x�����6>	;�cYX�S,od�HK�0�i��ᓎ���o�m�Z/�ӻO-f�U�F�c�7m�����	����;YXj�̓(�$���H17���x�ӻG�.��Y_y�vv�	�tww���mrTRFq�+ι��nY�tj�?Ŗ���uY�{砑y�o��6�1��"��5�7#��1Yʴ�	��ϙL�x��+Q��&+��Z���Y�=�3�֖q�K]�*:I�����$!���t�Z(q�oXI�jdB]t�0 "ÛKΊQ߅��	jɐ�>�!Tz���}b�d)�`3�]��m�Łs\��=��=��e��m슧ў�  ��vM��*�Jҧ���'C�y\F��F�*?r9;�uM��I -v��R?Zy�">�IY�s�ʍR�=�-A�<�?ݓ���)�P��vX����{��1x̤j��Z�c&��O��{�j ��c>�4wp����Db�w]~��"�;j4�^��r7W���t:�0@����;y�o�/�xzX«��J�3b�v?�
��Q�^n���8��8  �y作���5H�TT��\U��XNym�3�����k~��ƏwC��J�H�Ny����|�l᪑)�=����'V������ ��^7cI�ǧ#[e��̜�O���!98p� ���欕�`eF��E�Y��z���b7�(�)���1Ż������ԥ�~4�� ��$21{P�[��_=��V_8�������%����#
����b�����3?��.�Ow@�^���H��t�޶��/L
dW���_��I�:��J�.pG�}��`�eQ~3>�/��A���:Y9��a��5q�Lpr��;&U�a�6*����.����a.C	��u�ջ"$3"0�2F Y(.R�^*��;��+�E�h�|��7϶��]-��\y5Iư,O��2F5���"oڶ����P�/����=Ah>�j%��9��
ճ�����T�����C1�31�w����L!�����
l�ɚ&��s��c����R��D�<RS��:�wc������W}�Z�ꊲ�ȁ��>���T���1_�~�w�Db��޹A�v!<TA�,^<E��BF�>ZX5�k�~Cd�Y$�
wÎs
f��&��@v���v��s�� �:�+�Β��,��yw�5�xr��G�a*+.�pZ:�B��/�?"��Ⱥ�F�ۋI�,���xs(�0_J�v��;W�3w�-Y��\����������Opr�Ao����5�čM+�ѯ׵�P�^�i|�puc��VϪ� gd���������-�9��ɗU��0|Co+�b�o�2Avn��ʱ�H�$p���5�w?Ұ�����+�
%3�B�q\i�>�8�@��ꒈ�q��G�N�sYA��5�(�"�Hy��l��Dc������9�b����>b&fT��Ȧ2�C �(��g�	�
%�$�襒��QU��Sد
���K[�a���p(2�gr1 (��z�=�9�Ш��&�H��D1�������-��(�".�ءF�� ˋ�و��S�W�P��������m��N����<u��Wu�x����H��S8D�܏�q�;f6�4�v��հ�uA��%�4%5H"���= y�1���������*����Eo\���uә����I�F4�"�#b�k���,��g�f6?�;U}�j{-�W�� /	�x�P�nĠ�
��n'�+���\J��OQ���q$"��$�S�J�8ƳD���C�. ~�o��$8F#��/r>󞆫�ſ�A��>E�~K�;���&����Q�ꛡ?hq_�~&s$�V��Y�|Q%u�i�B��hM0ۆ��"/Ɛ�O�'=��Եa�I����J�������e��%�ҀH���EM��,/S�?�D���O'�AO��g�h˔4�A�\����Y�b�:'͎����'Lc~�3^�D���G_�����$�v�OC��-�����?���@]"��J��<��A�����q�Ue)s	p�HbԽ��w>Wćf�/�u`�JA[w�o��u�����4�%�#�4�.�RJg�-\/��g�Q��{�|�gTN��[�)�
�MҫA�9	���c�W�zӎڽq'�E;HG01���-���+p{
6$����Wo�:��MF���fv��f�4»Őh!�s�g�A�p�IL���c-u�N�����)X'k�ȖYQ�N����7������7��B���R0z��	�:�8F�o���ԕ�)��keO��ӱ�MV�S>po�/M�J��mJ	(U�ӎi�V�A P�N_i{ �H!A����s�;ć_t<!��ƥJ�3��_.�$����E��:����s>�S��<��+��)�/Ma��{qX�1���e���ڧ��G���.S�>&j"��~[�´L��onYu�n˺SG�0����jG_����+��#����ی��N��t�9����X����k���g�ĳU�we,�ڥ��tM�ӾV�{;+ks`�h�K	?��[�U"u��#| z>6m�}��z�]������)��ltĉ�O��I+t\ac&_W���4��-U/cO�pܜ��U���J��ݸog#=��s�Bh-�(�TyuyS�@��{����BES�l0�9OBPqO�B?���5Kh�n�3��B��Ry���ѴX	�
/���w�VB��"��SY�e���t�8'�UG�I��W
ζ��H������#v%3*�k}n�coO�j�g�*ptTN��"n,�W4_��;bª80������[�D\�$�:��Q0����S w"i�x������]������X�-um �}Ko�P�b7�~�3QY6U���P�z��R����<�U� �)\/K��w�L[}1A��9JM����y����=3������_,�[�#�w�Lm��H�wEiV�8W^	;�2�ն�GN臚f��a�>��(چ	�������'���r��~��I?++����<K>j���O�B}iW&�ڶo)$�|�4�۩�;Š)dc�!�j}�vs����W�U2�=܋$ooL��4��+TΡ,݇eC���|Į�:k�5�I�?���Q��o�� ��ٯi�������g�u�&��՝���cL4���{ն��.n��Z�P�䉨�$�P��vzK�r�D�%��U�f�=�Ps�~0H�?�ԙY�����Ȝ>��#|nh3u)�'u\ד3lr̽��g�n�Z~k� �mrXWtߤg�0�xH�z�w;�7)�+ pIJ��: �e�ypG��޽OI׫�H�\(�'���Ua�S9L����] ��J�o@��
]'��ꊆ��Ǐ�b-D9��~�)
쯝!�D�XM�o�����`o� �b_K�_��=�������NQ/�ڰ��ķ�T*�WS�0�s� |@���Q��T�kTJ�$Tcq�?�����=����S9�Z]�[Ə�����?q�.�%����?�Dwǎ�裏&#�p�F�(_Ck֖R�����9ulv>?��Dh�J*�ї��VBy��>8k��2�N�|���5sf�|���>ӊ�U�.�� >f�u�LW^y9u�O3N��2�F| �"5�a�z��gì7H55u��2������?�T���/���������C�a��.����A��.a�ʕ�F�U����w�Ü�
t�Q���ߓ���./��t�J���~��ʶ�;s?�0d�զA���=���1*�#�1�
�����i(p����������ߗ�)e��c��~�q*-]Cy>����0��Ր�)�z�L�8�y�B���T�R��ǐ��<p5)�*���i��/����P߾}��4z��_��W<�x���P���V]�VZ�t%�0 w�o}M	D3��`fa��ul�[_���<�\�p�$����@�^�CѰJ#��B��Q��������~���|�̥р�}��%ũ���f�z��<��^�֮[Eu5���ϟO�7m���uDF-/�D�FO��/���n]����x�*����Abp|>8v�}�������$(���|p�Y����}��E�6��үi�UL[yL/��w�U�6��y�Q$lq�#p��}z�,Rn����䂿��Rԃ/�U�v��m�/嬟�d-� 6e%b��E�ԱS<�
��x+u�`�r��d�9_�IlH���?�<��xz	�q�i�����oyQ@>T��.@\ȁ	��W]u;s�>7��i�TX؅/YĻ$�#%+��d�jJZ^ڶ��:u)�+����� m޴�����iM��j��ch�"|��5k֌��%%	�*/���ϙ	����M�\{���*]J��EG~F�֮-�Ꚑ]l9@U�:*[W�Lⴶ���4�P�+;Ā���9�1 ��G ���'��'�� �����6��;Z��m��+)T���nZK�C����p�x�h��-4w�����A�!CQ�>�U������j���z���?����W��Fz�����30(���ѣa�E�xS80�z|A2<�o��CǮ�.�3y��(�08�4=L��,�mٲ�����8�^�o�2oPC���1�%�/�0��0 ��\D��y�ƏF�:���ҕ|m���(&-_��j됴.E��A���N��������իv�m]�w N��JQ����W��9�|n޴�^{�E:��)�>Y�a-{ư!(�e�__���	�-���#���C�zı���]���.��
P���JgMǃ���Ac�r�F�֮YF��WR,VE>R�&ȃt��o�<o���~D�5	��۱�0�#0aT4���j�.��K=�#����?�����G���V��+nG��䥗�kdz�s�"�t�T[g�דφU[Q��8�$�[n���)�{��٠[YY�.\��Q�F��(���о�m]t�>˖|I��7?[�N�hU�reo���D�)Z���o;ڴ1D	�K7�p+���y�>���|��t�L?�}l�#p�WΙ9�QW�Ϡ}�G�z�^}�?�����)�{��tđ�r����5�LD�A�QUU-���@���ʫh�I� h�>�(h�6<�r�<��s,y�a��T�38��sU,AL��+3n A^���i$��IR<
�~,~���h���޼�i{e�?����O�K��u�_�=�Ye.@q�Yԛ�C���#x�k��o��ϋ��a;�@:��Q�1��ø��&�
GԾ}7�2�H�D=���6�����2k�!ھ}���;��4v�g�}�����w� u�������|����u�d]s�5�[زq=�{�%<�7u+�H�W,���6;�;*�%h�7�(�C�_������^�3N��y�OӺ5k�8�����r��!�Z?�Pv.��%]L�J����?��:��R�n;U�l�bҜ���i�hݺ
*��Fյ�}ޅ����{���w����d�>x�W^y��}��!0����@rA��u����LI�C��6�	~�@�$D�'�Q�C�(C�> ���K��oSUu��� !=:\���7�J$��������i�?�۴v��'N؟ƌ:H��'b�1�<�����d�Cy��dz�9:���q��H��g猷�z+��C�5ft������4�#���nc��*�B���4�d"BK����D-�UUo�H���>�c	2� ���Bk�ld�m�Y���I��'�y��ѳ�=G���6� ��Fh�$ZG��O��舩G�9g�I5U���I2'�u�z�Ek(/_��HY^
��Q����P^�*9�l�!�4�����p}��]v�et�����T^^��@;�� " ��. �C܋#�2�[층C��WD
zUvB����:� =OЖ���ʸ�����S�~�bfgVt�_�>�Y�q��i��8��<�ݾ��:w�gy�5T1o@����H$T1x�l�k�Oe��y�*� �:�;�<*�ѝz�!��1���#/8}`�=��C.L��O<��:�(���5�T^V��!�����C��C�E/-Y���7�8�|ew�i���胏?�pK��>�x�6��7��ɼQ<�d�w��t�Yg�AÆP,RK�U[��r��8"Q+�d�^Г0�F��H�G�������/���x 9^��	��#!�����R��X���D����M�雯>���j
�}*7�O���─px|D^?8��L���c��/W�w�t_��8`��7�?%���[����U�D�Y!Ês�GdL�rN/x���ٷ� α��T��OU�CN}�ʉ9��g_PM5损~��0�í;|�P'��|0���do���v��`��F�j�����G��W�i�F�rĀM6�~��!�P��9�D����#�������z�x���4���l�>`�lauG�M�<�N;�T�ٳ;��VQ2���3G������CAC8�î۷��	�@�g�[(��u xб#�� T]�u��JE/|�����2�2В�g���i���H�8}-��y��L��iS����T����={��h���>�d�@8)�'ڎ�$H�I�'6��Y�(��2qm��R�Cg$�|�53i�hX�6�PR{�N���R�G���<<�˚�W�ʕ��r]�̰XK��
l�f<�D�Ka�+m�}%�0�2&^)�g��� ��&��NU��ţ!WOD� n��#*�ߏ$��j:��{��, &g�M ��eRׂB:��cXY�=��Gh^)hc�n������!�O;�:u*u�܁�-�џ��L��s���^�U�V����`�׏��Z�1���i᢯�w��[���1��T �G��:��?�A,���S�$vk����*C�eu��WL�,��փ����C��q��m�����x[��o� F�!���oLd�|����|�s޹��c�q�8 �A0 J&����^ �-^�m߾�>s��d\mg�yLQ���@ｿ��a$*A�i���z��co����D{x�n���[��7��&/��A[�L}�	���:�Sg� Ε8e�Ef�.y�)�+I�dao0�C�����p�ް�����"�8O���[{ђ�幄�D�ޭ �,��G�^Y�2�������	��l#3J�F����R; ���<d�a�MR^~'�<�p�/Š(�|\���\1̲8h�w��s�,��j�5���!+�|�|��ǻ�5d�`���0)�>E��	�1�H�_,`�eH�P�����4�7��G��)� �	w�ѣG�ĉӞ8�M�3�H�~�U�Ѕ�ϋ��%D"|=p}��G��(�+��������.��w���3�������z&h��iC�J%��1�DurMP?y�v�F�;�S��Kp��xRe�D\��bٚ�����Y`c����r_�/�#�s�^��8�3W|'Z����8�8Ydd!�׽+�,���@�%ͷ$��;��v�eW�FԂ'�+�"���) �c��[v���󥾄 ��&� iJ�E@[ȿԻ@_�x����kQ�I�O�w�}��_J>3E�D2�>#)�� %y����Qu�h;�б�<� ��GT��~��ڸ��~w�oc+�?��G��]��c��ǜ9s�D��_"��%0����!�"E�eG�>GL�E�@�{,ؒ.�	��
������vR"w�ഖ�6����$��a0 �m�F� gܸ���v���D͐ÿ�b��z+}�����/2^���g��#G�y�����Z��cၫ'4�>"�ҧioJQ�f;��B�(�f?�R���������>��:�*����ۧ��L�j�}t�Z�P�|�  �F.�s�'1r�}��/@+�X��~�i�jc�$x�#�
-����E��sJ2.NyN]C籱�H�~�|J�|�� ��� ���Y}7%�,��]zۤo�|��ޘ빂�|?�To��c���CGR
	�L"V� �RA��ku�\@E�=9
�5}�"N��r���!��&v����O�;�z ����pA�0�y睼c�Dh3�;�v��(�`d�1[�h>X� �ʐ���?\XTpe��i%�������a�hDe~T@Z�dᓉ*�������<0T&����@�2R�"�
�P���q�����s��>���O*߾��"���@����j�"ڼ���*D�f�Fzo�'�d�챐��Ճ���k���K�]c�	}&�4�
`�J&�l�dLu�_^�e�B�H�Ut@����:��6�_�r�����
l��,$2�B�0�E��.� Y�t�^��m���N�Rr�>)D$�+�Q��Y(	}.I���`G����+�0hp�	����G�+���@G�7pu+�G^�H!/��F�n�����;v�	����{��x�ͷ�G�|���#.�����v����(ʉ,��C��O�%d ���� �%��HLͿ�c�\�^�I&\&���ŕ�`�֪��)��,&%2�q����ė��q�G�|��CI�!�i��G�d��8�A2RaZ�v)�Z��k��^Z�v͝�1��*�����5�\ku�d��'ͽ+%� @���g�E ����`ӵ^L^	�G_bl�ѩI�����'=d_
wX�s�w𿠦p}�nF�`<ڀk�}E9�3
 $���e"�c�w�L�_��SG��<�h�����˞���~�/���P�}w����x�V1�Ȅ�X��=���~4��IdQs!Y[�s�X�9p�>���y�F�����@�����[hђ��������@�z!�3(]��t-� n������@d�q�$�t�v?��

��5k��m��9mz��U���f��(���D��\�.����f��Ź�q��`�|�ǵ�L��~�v �>Ĉ�E��^����P���6Њe_S<���@�JK7л�>J�����r�	�plk<��L��"�Z�k�a��h��������ݔ�1������ୁ������v2V� }�<� ��y�E�Ƃ$;H</�{8�%���0�b?��1��)���� &;F�%��*#��L��DD)<��(4rd;O(h3�Aa��]��c��㑘���a�d�v E>�z�J�HE��&��7n�rD���C&<�z�N�(�x�����|ҢD
6b��kp,j���+�p�1��9�}�)]����B�!��E��cA�� :�J�CY�kd�(��nW��1.���"�4�6��5|ݧq��G��k�2x�Q�V_���߲ʋ�&a��	m� �#x?�t��P�����~���?L7�����Q�I(Բn�&zw�'\��4����O��;x��V�G; ~�?�8�O�X���� _{��B�SO=œOvm22Q��Ȯ�>F�$�ɵtZ�Q{�^` Zl��Q�M]�������N���0��er�f'FTD}��w~>����4�u0?�s�[ ��믳���_b��/�g���}�a�~��/~� Bd����K�&��v�(ϔ�=� 8j�6�#����H��b��b�^����P"�����JZ0b�TVM.�J���y~���p+J����g��;{�%R<�.��5�,��GqE����x�]�Г���c�1 S��w��߲����;���`3�ْ��)�.���	��B&���̚� &2���|:_=G�(��|/m�\F>���&����B0ОV�*�y|F�*�컌�?}���&��ښ��<s�L�P�\QO^�LLq)6��	��l��0�Ђ�r����x��y�B mF7,$�uY��#*Z��a�9��LP�"`�äǳ~���gM���y�~�I�&�_D��,���]`����{Pp.�{�M��rr,vx6��xθ&+ v�9�ոq��Ya��������B�+�'��Xu���h��)%�{1���t��jN�fQ2UG�L�'�"�7��OI��ӀA#�������@�s�@6�r?��@�讶>�M<v��s�����D���:N	���j�Yz`ZI�_C�ʋ��>lԁU�vݒ�!��354���y.@9��|�h����w)���D˗~�Y=M�Q���Z���U������k��b1(�8���j�hъ�m}��7�A�`Q���1�-0��Ȑ�K.I�'�Z�,��t(��Ď��������f`��O~����#�0��?b ���3�h x}�_Z!*���\W�S*Z�Î�B�Wp���N`� 9�v�L���n�İ8��x1DPǊh��B9��7�a����]w/��=��=�=�-���P�K�����1���$vK$�h��h"�t�㬷�t��`�R��]8���A���ߟg�tFb7esB�8�9��͝�믲3���z&;  �k�uA0E�[l��ؤ�z�����'m��w�2�]�a�.�������$��t�]u:(� �3�Mhcp	e��j�	Z�b1��[N>�E~o��Q���'��|;���TFY���Ę�4�?s��=�@h��U� S��16���x�@� 8A�������>~�\�VB��K/����cq.���(�@��Y���������_.��_q��)������}�g����TԮh�h@���{���
��BH�,B(����X�d�õ�;Eܐ+�`��n �� �yj�̺�)�@�����Z�\�?���v�x��<i,E�8�c�R�&�׿.gWϣ�:���	�n��~C1�_�{����>����_BpAD��E3�>�3ĉ��XY�Equ��
�~2g��'2��9|�%G�\�	�E��#����%�.=�K��m�����Ȁ6�����	��@�d���b$h��o(T�|��f���]!���\����y�C����O$�5�N %�֚iDO#H�4*�q�k;���KJ� $�;$�B�t�E�@��?!�4=?��#�W>��w��~;����?�1�eq�<�{�w HaW�����ڴi������T���x ��1�(&LH{��>�"�	�h<�	8���L9�98��-�]���s.B.�+D���u`�s�y���E�w4���!�0vM�:�,� ���
�t���	\u���'R4nq�^s����#�3(�?�r��������8�]z]��y���ϐaQ:uW�F4�p�iO�BU�d�}t#��ً6���� ����x��; '~YY~��;�` ��Zj�o�����27    IDAT�(���ƊFԾC7Z_���.+��0"|���߷O۝�u�t�xa ��I18
� @��M��c)�iUF�����uA�����y��ǩg�^�9#�hZ�׿���TPX��x�hh��^�S���c�� ȣ��,V��@����5cG��K ��\�7���6j�Е��5���of�4Y�s�-C�c�wh��E`����i��c��;�B"FmQ��ZN�;~��zVO��f���NЏLJ�$bI�s�.��#�Q )C��<^������b0�/]�2c//ڤ�� �sYGd|:G����~N�aQ��g??��mP�o����P=bm��
t�1�g癑�Y���89'�^U�ro�l����-j�b�0����!�9H��Q�<������˧X"ɉ��O={(͂�����Ř�P
�/솤��h�H�'5@р�����c� ��9@������y�^��c���`���7���� p�\�]Py�߇~�;�@
P�1c�a! �ʽ8��&�馛ҁ� g|�Pa�B�kKIP^Ai�3��#�7d�G���>��)Y$|C6�},hX\�N�+�K���E��}�$^�I�w�﹂��硔!���R��ԑ��d��~��?Ծ]g6�r��]��J��rTSU���s�EC�|�wI:8Ѿ�0"�� �3[�n�'��􀓟�l�d��X(L(�x�`� `�K�-�X�w�q�_�^�8�'&�cnJ�ʕ�i�ܷ�&���~���~;�Y=��mՒϛ��%܏z�(TG��Z/�Ȑ�H�J�ᢿ�cE;�/���>c��!T�ѷX�la=x�Hv�D�\ �C�@Rn�H������q<�����������<�'�P��*<_Q>����Ba1B;�o_\[E�p/����!��RAN�y�� Ա�by�[�v�W_}�89_vI�����F��kz'����sp��D-u��P���k)�qv[D�#�-�z"���ǞH�����s����<~P�w���ڎ�$��9��f��3;�Ocm�!�9�W��u�7I�늑�@��ud�\=ۮ�C��l�d[��~�cF��ɇM��p��l��2�!�xSL	��N��|ݗW�� b��DRɫ�k�Sgٲo��l5�=d%c�1*H�={��\]A�|�5UVE8�F���Ѐ��Ͽ�k����q � ��N:��W=�I4T�%:�b��X4` �5j11ax=�i���L�`��w5vH&���ջ7�
 ��~���.���i��;���ޡEc\Q����y�B������d`�Q]����?��ϋk'vH���(hY���C&���}�;p�0�"�0��XH$L��+�
	@�	H�*�7�<�&����)i�q��.�\V�*e/+�ѣ�҄	�ϓ�?�����~�~k�}ߗtB����� #�ҝaT@@ �E��8��1&�0Bt=���â��d�I��{-�W�V뭻��|���[��Mխ�y[��=�Ou������<���<�͟��T��FƊ6o�b�����X���I2�����=wr"�ց7Y���D,��zW���;�|���^�}_(��yԺ{{�g$Pd(��e�d�+�V�#&)zF<�����k^�j��h��3aae��3�Kֈ��8R鏍��:`���W���F(�`<=�i~29��F��UO�!T�x�N�d�h�\���(|3��Z�r��{�x��6R�K:���z�+(�E���qu���(a��r84�g���\t��y`>_�!��0G6Z�={\�%��G�eB���#�g������B���8�	��^�{�ġ��ݻ����QQ�0i���c��*<'J��SJ
�;4yNA�%��,�Q�<��r���;&B=�p�"dyw| r�J��u���p��5�o �չ��g�^�5�������`==��÷^�͛�{y�L��Ț�綶�V��P�YG�l���W�x��{9���fQ�4{
�~�w��<31/�(>Y��}2���ԟ�w��VB�5�f�:W*�-[�,�xa��T��*���l�����s{)�R���)�q3�f�@,�f������wO��'">���k�m"���m[��*L����X�`�KkU�c�a6/�	�S,�ȨdQ=���D�;^�[�z�N��ju��Y�~��^-Z�����y�sx����6:V�F�bfk׭��+����]ҙM��I�}��#"'\�C?���f2��į����#�F��ɣ�C���@D4��v]�M�0�c����;~��qo�q��C�&@
 ��ً�Z@])E�KX�S�XZ��}Շ�"�uP���(�1��@����n��5{�!͟5��A�4Ԑ�p3���<�G���z���|&a��y۹�^�-�(Y:Y��n��Z��iu�9���q��24Hi�X!����Ü������uA�l,s�k��f�w(a�;�B�e��((���n��;za�cHpO��:���6�4��������mOJ�6��ͥ�^��/���0]3%h�yX�t�z�+��>�D�N�:a<�]ג\���m���U��\�ȑv7á&��DGH��h��Ֆ����p|��Oʢ������n;3�P��\�;��2���}���6:ְF*��TճQ'R�Ǘ�T�̉F�ɘ�zPYߠq�b��`s6������Fи�����/|�A�Z��U>�s�\���ż��������)@���8v�r]���'��7�r�SWh��L����G�#�'a҇
QE�P*�wı�D;()KB�{f�S��¢�^��L�?Z+q�X�X���c�<����>���͋��7_w��_��V�^i54Vr*u�ow�g����~���y���˦)�@?�e��{������b��ɢ��p�ʅ!��S��#���ظ��x�����v�?|�P~��2Q���?�8͙�e�LچG��g����M��K��ƍW��;<�R��U��̳OM�8	:l��z�>�5���w*�_�4k��K읿�v��l�T�a}G{o�J�d�Lڵ���CL[�i�������y\ D� �4
�cҵQ �"I����w���hf����<9筷�;u�ی��H���;`8���q`�[�Ɩ/���|�����7��K^k��y]�	�Xiˊ�bnЖѬ���7�D�G;&��_ו������	�����?����^����-�ͺ����l��:d��r\�[
�h�0��A(.c�x@|�3���'����J
��p��1�x������c	��@���IL�
�M���� ?�O�u�[V��T3���<q�>���5sI%�Z��nW��F/�ݺuvͳ��|�l���dl%��C�8ξ��x~���?��I����eng��f�XC�x�T@ɲc~8�d�ŋ8M{��I{��'m�L��ǜV�g۬X�x�E�����l��%�\����V�Xa�Q�X���i�={�xhh�����dO|��׿��v�O]���~;u�=�k�ϟ�S'�˲�H�ldp���Z笥����c�S�cO��dN���N1�_~4�OZ���:�)�3���#g-�L[&�a==��U��86��&������ݏ-�Ϙ@��1�R��B�㌖̢��������LlEca��b9��7{��; �X�YE-���͋�G��x�?�2�gh�>�`��gº����7���;o������ODٽ�i�7k�����)18�y^����ONe'#9�6 �� �!G�
����B�`)�
�F� ��/��K��M��ۮ�-�iX�D+G�ի7ؚ��Xjxm�l6�a�����yFm���(l�&Nw��F�}"m��G졇�^����J@맪't��uyn�
�U�kTG��w�����J�UR�V-��[�a6^(��c�v����7���$��_��_��u�Ȣf�'.�v�����/6��O|���=�������&����Ä��}���|�b�U��o��/m붫lt����?�ٰ,5AJ劝<~ʆF+6p�lo��o�9@�Z99O�c�������R�?��Y�<f�d�Μ9b�=k��l��Y��?mc�����������㣈*7���`��%rg��s P6'��E3f�J�D��QCu�K��ht<�?�g���#��2��ٖ�[=�h�O�s��#��ޫp�2��١c�����J�'|O��BOhМ�c�	*JH�� @IF���}�"@H�C  ����]@(@��	T��8��|��O*Y��������K�Imݚ�m���,���*�`=_B8�;:]��5�8|Q* ��z�(��o}���X;U�|G()��k��<��J���=k�ʈ5�e�;�g��H,sK2�fǏ��b�aǎ�[��N۾�j��=��<H�G��d�ό�[���������J��{����ۿ�V�n�j�?�h�]���"���b1r �r����<6`��,;|d�6l��)Z%� ڀI��Y3�ACCӜULG��^�÷2^���\�a=={���V#q(�m��� �i�B�2�>�l��e�F�9��h�܌;>8ru�b���,B�(@���d�Q=�lp�)�+ |��;��/��"��=�:B�G����@�a]P3�?4�# �5Ƚ h-B1�.��8�cD9�
e��\�*�rh�q�����p�N���`9p}�'h�XXD�`A�(�(i��fM��B����i��E�D����\�m�Ԯ޵���%��m�u�Zd�_q�Y��J���HeL��'�X�Fl|�>���@1����o���Zd��Ԕ"� _!����c8~h�����l�ڥN=��+ǭ���}
�Z���=쾉ѱ��Z�����wXG�l;yj��z��S��[v�ghx�C�4Қ�+�W?�^/��ݳ���7��y�c�{�4N(5M�mhpغ�{�����c[�&�I�X���h�T=#��DLl68q�ԅ<�ٜ���p���IT=sq�8lgN���[+�[ �筯�k�����sV_ �_�3o��4'8{���Q�)�q%�B�=�*����P. ��������誉
�g� ��C�q�j�ε8O�;�& .JJ�E�9�/�%�&��r�u��T�kI �x�St���C�����uT��5۸����|3��KY�e\�#
�$,a�PO�8��������_*[.�r�/��յҮܴ�2�v��	�C@5��8~|rQ����sv�0A�1��94|�֔2���r�X "ð��������|�6o�`����w����b���B�n�=w�2��v��/7�S�|�
��7R����۩��x����u�݃�C�>��=�6�j����T�f���}��u����^�����6>Vp��d�l���9r�R�Y����bӎ	�gS�� W����H�4�8�S�Ntc�l�yq����D�j'���=�X�FB���Ȓ = ���z���J���X�("�y15-�8z��[�x�d2���_߻�4Τ�,��TV�����k�������Щ�s���y�����M��Rք�		��1���ֈ�wx|�<�YϦ���u�q�[���Tb�����*߅��`_�g:���/Xow�����l��Wx��<�u������k�o���h�r۵�Z��Ky�Wwx{;Ԇ�������D� ������U�ư�H�D��̄�B��88�}��_�(�9sf��C�}L�wTm߾nK����Q+V������jG�#�K�qԺ����En���}�|bhh�7��=&���������w��_����~�N8}�J�b�O��P,ّ��66^���5��ҫܳ���I6�q��MQl/�+���(,���*��'~�^�h��>���O=lgΞ�������:M�H[6�n}GO۷�����,��l���d�ǛX\<�o3� (�T���&i��p	����څ]\"A�^��N�y�ֵqB�-v�K�I�&���h�uX��.V�tr��}	E�85F�v���,l���8��^=ח�YA�r��zg:p��y���m�%�b���'�k���C͈���ވ���uA���n	+Z�Z�(�T��͌U�)�5�~��W[��o�6+�	���x\����#�4�^4���}L�oYc8�J×D>�|'�D�#�����)����b��-����?y̪��[��2/�O&�e�N���K���?d��s���1�����+�_�p��fjI����gQΞ�i�|��l��%�ޖ���_�+�Z�6�_L?�;��Œ�����Ƭ�t����w�㌍I�6&E����LD �S�� ���jT�W+��h�,sm�<qB�9`'Ou��\)xUO�Rx/��}z�>i��,7:�f�r��?tBJR���M���P|����Pb!�zC�V@h;��&�^Cm\�ǉ+�Ix~��f�s��4��u�P#��s����9�/IJ���P�,�����	�PP��-�f�L�j(�4�\;l��K��b��Y�{����3~��8�{����|.e�zɮ�b��ܹ�s`���wȵ�{M���k	[�z�U=�&�}/��I|��>g��/����;��N{�k~ƅyDt1O�����N��O��r�>��}�ha��S	;5pʊ�1�1� �z����q������7~�k](}��G=˻T�|�/��$���w����Ї'���j%�F�[n�����6V�F�h���sV��G!X4s��e��6tn�N��5Kvٛ�����<B�T��E ȓ~Ы�
�:�Y({���I$B�	gQ���*�P��>Lzil�Ν;c�:����Y:8�̒�W��И������k����k�y�8�E�}BS?����� �ٔ5GY��k~*�����E�7�����e�:�����t�/KA>	���-�
QNa$����)ԶC�Z,�@W���JX{du�,�4���JP7[*/U�!�/��kVZ�&�?��7��O9�R�9]Y�;���uG�xT�����Ȗ�x�t�KĹ�X |::���@�D��������O��!��R����������ر�����;2|�
�v�d���7Jʹ��:�y�IK����s{�E�?�V[�d������w����po�
b�^�ɝ�n�����M	���Ă^�|���]�b�ͷbaԆG��#�|����D#2)�eʽ���c��̳k����L2�rl Ջ�!�VzQ�S<p�lZ8B��r�h���6�&����5��g��=K'1�Փ��|QS�0�k��B�H�Y�v�z3��	���"!.�� ���7���4�f�#&ː��<iѡ�>ḇ�G ;-���}�Ly����.��9�C/C�<�eB���Ofq�<�q�Ӹ���BJ(����T�<%��f�n�g�Q�����-�({�Wi|��u5�Q�e"��b�b�sl��^�'s���p$����V-����)��p�b1�Z���C6:%�(#��(!�����[�*6p��>t�N�������6K4�^_��Jf슍[l��U^���@�,�p�M6v�Fc��h�x��TEB\�u�ַ���Fm��.;sf���N�BR�}�Nۺ}�D��K�B���u�?� p|�m���P/��<0�	�ęL($Rǽ�b*��'�}�8���Þ^�j�ly��b��6^�������M ��������{��Es�����oH?4[�=�/� i�D�6-�?3QP:Oc��!@���|�eYH��y�V��]�#��� Y�u��K��*,�&�3�4����v+������m����L����E�H@�X����,YBmh��F��XH�@�.��a����z�T��W�	��I�ܰ�J��[�yKPJ�����w�    IDATa�1�>0p�>��>g�Ҹ+R�Qf�*�K�w%��P���	�ݳ�+�
֖�X__�=���=4���âF�+V���o���̙��B�9��E9tz��gF��n������_�J�WU�Z��Y,�{ӊ��Fn���I;E�0o�Y���p����=���Q�(&���:���P%,TZ�7����T��@�ؖ���5m6ɲ 8@ǿ�~�N��X��=q{:�p���{���=f�c��f�^%��[�bu$$�+�x�>���GH��+c�����;�R���m�N%<D{|��K���t/Γ�PXg���<��s��9�<r�N��J
�yo�y�B���C��g���ZD )�?�~B�*O�
?�'�����][�P��7P��J�D��U��j�T#�?����Ջ�}�e��͖�G�I���w(������1��"�oo���>h�����y�����w� ����16�C�w�hb?��
7V�U��`���J�IgG�G���%'%0%�����xN�9h�o~���v,��%�Qѹ�>3�o�s���{%�D����.�ȭ[7{���~����{z�%HĿ>���.��nB�S-5�&,�E� `A�!J�Ϳ{��y�E�ڏ��T~tޟ�rq@�U���,۾��@�/�z�liZ?&���s��i���R�膜7���K�)�-.nIg9 
9cƀM�u���D?1��Y�*Q�xJ �2��/ R�fb��p"��P�G`c�q<�AT�^c����9��p׆� #ƞg&v���]�~d��X(�D�l5�x�,lz	M6� �g�W�%����[��{�X��D�����pMţ��Y��	���?W���M%
��g,�G�J��%ͼqnX�q$�AIz/]������	O�"ڇz��,А�y^}�&+Ǽ��$v5��'i�5{�]�e�G Q�n^hހ?-�3������w���ٟ?��M���\@��G���}����Ԍ��E����[}	%oԫ�k˻J��7�I%��D}��oG�qw�tTl���,����i��1������+lێ�v�����Ʉ�g�r`ч�t���A�%ٚ$uQ3���L���OD��6��#����[5s����#�m�T��k%��F-���B Q���}}�v���c�굤�]�>���{�.�CI[�j1�� �f �qz!`�v�V$)������a���G13	U�Yuo(�FF%�qŜ�: !ay��l<
�~+͘��l	��������͍�M���4�H ��zTڤ\��}�A�l\(��F.�$�OB��|��'�G�Y�Ō�Z6�.܃�PuX�EX�=nٲş�h
"@�*V$�+�'������Qh��'�źe�B?��Bk�8� Y`<Ϗ��5�j��U�P�0�{'�����&�.��	���Q=���m��N����^�皫7��)ژNd�TnX�m���3w�OC��:��6��j�Q����g����w�����n��V��#ܓcM�?B����߉R�>q�w���Q�Q@j'��")���ɧ��y@�Jd��]��'��L�󟺼CӨi@e�+CVC�c1���dܵxMJ=������I�' P��?�A��{|)S� �0Z�����j���9}�z?g�҈�57sm]v��xTۇ�΀������3/ry�K���j	���Q@���#��	�c��ËEŘQs���%@�	� 4(�����E�y��G�MŘ�`G���G  Ҙ�gxX
�Q����� U�m�|��ا?�ihr4e">���fF � P9���F+$������^]��C  Y�J�`� ̈�WD�.��@E��]��A�I,�Y#�1`iV����r8l��y#f��C�I�����Ġ&e#�;�G�ERm���<�04ɅX-���� ��$�"��*��9����g��zz[6ٰjm̶m��v��̊��FK-a�L���Zn�6l��IZ��Jw�jO�?<;�V�
��}�3 P1o{���C�kpg<QX(�G�&(�ЂcND)�*7�NtR@O�'�1�¨�h��o�u�g���?�#Gd���Z��u՛9_E�4K_-��-@`�g�e��� h��[����W�j�d]�.��������iTk^ҹ��ɉ�nQ3�FT������.3� '�ECcs��Y��� �G?�Q{�k^��-��L�� F�B[D@0/l@�z��Z�	Z�� 	@��Jm ��4rd����c4��kM�b�U���<� �l� �(�v-.B:g>@(����;k�͏@C�N�0@���Z@�G���'
�!T~4��ތ-��&H��d]!����ð`X�|�*���I_c��cҌ	sûBePH��5<7�KDy��"4��v�!�0@h�>܏�X�|Tj�#'���J:������@TϿ��r)�re�vn�ܶo��C����<.���XǬ�6>^�j\ٓ`	�ѕ�j9�ԫ^6����
���}�{<��g�b	a��֩�
�KM	X�5s�5��q�~���w�5�x�}Z,�j���XͿeU�x�B���P (��9�Z1�!'�̿q�����j���aΫQ�%�ܻ�����e��O����Nؓ������rVk�����#66vk��bY�����{�}������VҏLd�l��y�&
�r���D��� � ���1��$�Q�8x�cs"\��;�U?y>,1�h�9�ȓ���Ei�*;V����$n\��h� *-3P�� k �x���������]w�����@�g=�BQ	"@��L�6M�i����]ԑ�5� f���tPj\���E�	���L l�������a�b��bC��@�1N���xƇ���ȉ�����'̎n�W�6О]�$�����L\�?�ߊ����k��+��}�Wk�^j+�\i�:%*���4�N����LD�`&�t�A<V(x�^��GuPذ:��+S�RZ{�#��X(B4��/֏�����G2�5�[v�~Q�\����hIi�k���P�H�7��\
�G��;�1�, ���%��l��ג�M�^AC�ٹ���'�F�>�ԸOؑ�1��MN3��zRҙ���3�p����d��w��0XGP2l*U�d�Uvm ��PѪ��DB�;>|  ;�8�0�k3)���C@��riV�g��M-M�gCp��w�s�� �?��s"��]3��n���~Ο��������D���Y�\��P\��<��E�@��z��"� ��yg���̀���JQG_,,31��5�c�b�7��1�Z���`e�<ļ3�h�X#<��1Y9��J�\ɩ�B���������|�T;�k�F۾�rK����9��z�[��*�6�V�'�A��Z�����#~�<�b���r�|�9ғ���wG�S_|ƞ�fܨ.���|�~��0�K�-�I��!� ��hi����o1N����wF�����#��T!�#�r���Q6���ߘI�\hQ*��h��X
��h���k��7,�6;kǎ����yR�s����3�?�����������F� � ��)9 d��!�D�������C�x @�#xo��c��E�b̠'�ș b +� ;ԉ����� XC�\_�	�q�H�h68���������@��9~�"���t܃ka)��o�[����g�Fk�Fh��:2�� �j��
Nj��x���NW�AG��}�N�O�ϸpm			F���X.�(��@���c2�|x&(N,+Q��������&�d*Z�����q��1���*�^<����F�*6�R[�f�͞���;$29KT�zD�e,��ɦ]������>_�zT���c��T�9U�g�{	נhq�a��K�F0�\Kʢ"�Z�����n���}n�whh�=Sq�tih��Zf��t�Ĥ9M5��|Y ���hB�)'����A��7��ꓨZ�6j��!;s昝8�cV�!�_	�Kz��Ѩ���>4��G������@�KfY; �$�V\04`�JX�M7��9�GÇfPC�8�~E��^6��0�8�c�9�s�����8D���<#߳�)ԇ6�?�v��X�Zͩ�	x�ݰj��p�h�8����K�X��@ A�`=�}�4d=���7�e�@s�R �yg�1��yXT�3�$~���&4 ŸBc��2�9��	�*����!|��4R�C� �emx�z��~48q����2�p✃pVn��k̉O�S���9��Ba7���{���Q+�V����d�ƸY��c�,a��$;q��<���ͷy�;��h�T����;�z�h���P*<4�ֻ��Q�G�:o�@	;�£C�AX���J9l43W�e����{*�,���w�Tܿ��Pp��C�˹����5YD���s4$L~�^���0KT���G�T�eSu��j�&���NB=�����oT�?k��<� ������4PQ5
d18E����� Z'�1c�E�3�aB�) 8R����	x"Դ]4���
d���V���������w<�V�/4�k��b�p=��`m�vۻ��?BI B�{Q����Hy�6c�?�*�8[�l�J��G0����;����F���?A�T���gM3X<�/��cqM���r,ϧh"�Hh�r�ù�0h$�3��
���'��O3��[OOTҹn�y�Z����I��`Z&=�GJ6g�����a)��I���l��g\	#��λ��9ͷS!7:��yY�
"�~������؇�������l���-Xxیl�8�K�ntw�0�q�prB�j�2Y^2��[��8�l<b���h�o�bO?y�x�?qι4�a�nƶ��0���o����ڻl�P����g)�����S	.Z�DHP�Q22��R�o���3����^�"���dI�����cj-M��C�h��+sqmy9�B�D@������~���uq�P*PC�,��D!�y��XD� ����=Ѥ�%ᫌ�Ve�� �;��b�f�xVU��$r=��wFH��ܛkb0g֢��/���a�w#��5˹ⶹ&τ��傠��X��"��S!C���/њ��D�Oe��/Xo�a��?:v֮�z���S�l�0�;�L֪��n�:V�,���WY*M[Ժ��qͭ{�{��G�c��Oi��eh���B!�5�R�C�����R_g�
��֘07��ߕ��
[�y+����U`�s��ܥ}6[�'��,*�k��Z��1���N����A� �w����W-Q/��fuം�,�b%K1��ځ���Ǟ����'}���r����b5s�F�C�$�Yc	8C�����@���Q�ތ!�E�	�7��ax�"M�0И���$ņ|� ж�x�T�.�A̛�6�^f;@Z#<a|j̃���%�Z� �ϵe١y�
�û���������]є��.PK\ޝwCx�[ ��&?m+�֋�5�D�qo�K�1�r@h��:NYuSh��W�.�$j�ga�3P]�{��	�����Ԯ����=�MĚ�y�5� Z�w�*��^�vݼ�&8��+⪞�"9|)��qGj���M�m��+,��z�o�ޒtK���Za�dU/�\�|[�;~=�2���pl�+|��&ٓ<���\�Q�F�	�sQcr��]�5\g���p�$E�_�F�Z���,\����җ��������i��3�,X����Z�)TO&1�b�i*�xX��X��o�y�%幷��l��Bi6�j���h��IFo٪%
WQ�6�`_�elp�`�D�ʕ�,q�˗-�����0�a.tލ�6?!��s -�b��@	`@q��Frt�'����� T�7 e�����+�G<`�#�EH	\4�2�����hL9^��O���1�z�C[���%�U���yމw D�l~�#�����>Pp�D��`�6M�)`������P.��揟 ��Z�̬]�%|%aƅq@�p<�
M�{a����0��<B�s�P�^�R���A�u�_~Q'-@��\<�g�
/�|��D��Mٓ��kE��H��Ymf����)����@�'V�&��HY���\�͊�(@�8>�}F%�P�%ӕ����(2֒
���Pȅ�(�kM��0��f�*��Y����o��o�����ӄzJ"��*�]��f`s�  �]Z�jvȡ�w �4���S�!�P�tp�:F�)a�`���CV),�m�yu�(EͿTI�h�j����3:-_F���.nw9
%д	xW���`C! T�5 ��ln~'�@�)��#��i�r�|4t�08�*<6�~� x.�A~��&����>D�i��W+B-\�7�E�p}�(izh��MJ�뉱A;�U�F�O<�:�j�+34
�B!��/��%�9Z������� 0��DQpO��\0'�cM2����X�#Qb��S~"�p8�ySY
���r�<>#�V Z��h.�d� �~X4��XOO�u�wX�4b�d��U�4<J[��h���g�Ξ��6n�f	�zE���1��eU/��"n�駟}��|ܰڇg�0�����1d����h3�Z�̍���a����1dO�\�l�߳珇�o���+�����ĝ�Q�d^n�^���t%"�́F��l��
ȧ�Ρ���-\2��*ɋ�'��������Z��Z�D լAU�l����g��R#�n�/Yk+�/���HR��q�Ffч�Ei��5#�_��4om
EN��F����Fi�:�ߡ(�#E\pOi[�V�����

-/��d��y|�dѦ���ϵ���s�4QMat����QD��$�Bk��d���T�A��,S���hL�!ϫ,w���3+��Q��9��q_�%��k��Ƶ5��;O�o.�����cL�8�S���s˹�(چu���K�X�:�e��(y��i��;��x�n�V�}��N_�"h�h|3n�}�'#|h4\@Wc+k�C��;�
�C9\�1W=)�%�f�0D`C���A("4�(7~�20�OD{
���Ok���f0����%����:�� *�y4=8LņK L�
56�xa��{�c!���I&jv��S6����esIKԫ��ʣ-:���}灇md���x������5��bT�x்.��ؠŰ��=���yKi�l,�IZNH�79w%�Gi�y���X���ϩ�' �Uǵ��#%ABBڜ�Eq�l��tM"kI� DJ�~���7O���Z���9�g���y<oi��IWֹ�+t�A�r@r��Y'��X1ךC�'Q������ʟZ�Mt��:]�l&a�ڸ��v��tnT"���m�7��-�=�����:w�9��Yq�lt�i�Ko��;~�-���7�4AI���� 1���"k�c�
&V"V��=QG�&(�'(B�>�Kx%`*v�e�o��3	�+76��8��Xf��&4�"M�c�˄�z��8��H��{Q"'ؼd�NI�$��w�#6<|��U4\VQ�p����a����~�
cKg��J8��{��b���N�"�i�r�3C8��j৸T��j�(|�kl�fB�I�� �����p=6����k���mq���G�&��E �@��8_Z��$��>�X��:N�������B@E��}��r_{�IK0!Ƞĸ�4x����(���}=C(�$����$���CKq* �{Pҹ^����aˤ���!�r�z۹�*K6"��)�\�P��l��e�e�.+V�6,��{�&���F�-�?���>h���֬��N�=e������C �J�#c�>Ƿ���^�Z��QLQ4�����/�����>��>�B�>7���v㍯�&<I)�aw>���޼����_h[�l��wy��5�IDy`�� e*����A��c( �*ԓ�t�3v��a;}����/    IDATU�c���(���\~����?e�Σ�Б)�&��K�{}.V��(i���%8F��%zi�i��t!�0�3��K�4���e���I[�!(�u�*�%���s�kB�c�f,����OBCt����9*�gܸ�'�{*��"ǤK��K )�M�U�c��)�� ��Ѹs=	EJ5BY`�B~ 	E�I��&�?/ ������D�oV�M�а7Z&E�fT\.��]�,�d�lպKl���f��&b��'
�������OM�d(�K��d,�ې�Cd��Y��ɾｷ[[[��mY/�|��q{�{߷����o`Ū��;���a�t���Pw�����o�/h�/�����S��K�w���p�l�D�������Ν0h��� �U��⥫�k^i��Q�)�q�L��~E���ӂ���Q{<9�ظ�>��V��&�����f�L�Ϟ�Ç��b��k�C�g+9v���S���;ԓI^5����o^��¢;H��Zn��n|��@Z&?�'p�w�G�d�:�j����- ����F`���l��d�9N���Ӑ��=��7�D\O�o��hQ$�^xvmx	{i�>F��k~�ֈ�AE�	h$T[�~j���� ��.�z&���%�{zڧT�m[/��;6y���r�b�d�.{�.�5w�e3m��ztl�#���z�j5��l�C���Oz�s�LFY�a���5�ߎ+B]�Xw�2BUٕ+�Y�R�Ju�~���l���V��-�H�u��>�.�|�m�~��)A�L�����O#k�g �V��=����F�x	�¼��֭o��
�C66|�N���޽6Vt�ϻ��='�v����+I�;o����q��r�<�f$�[���Ą��O#
ca�
 Ĉ��*�� �Q:e����ؑ笧�+���\&c�|�uw������6�sA& ��F�L�A�����H��}fuF��DE���V�(c#�(cE�	ILQ��W�6E8'@U�i��[�7	ݛ���*��n���s ��Һe��9
r�[�{Y���k&�ώӏ1����y�$넱iV�uC��z���Um�����q�'r���m���M��b�F�/]mk.�ʒ�v+V�^�'�J{/���X�)K�纎2��Iu|�Ɍ;g�KE��z�����{���g���;�����ș�G��{�<�φG�hR��
R���F+���]��M��	+���hѾ�կ{QH��~�VY�/gny��J:k�9O�_�h���i��?��-Y:���<u��e4����ㅪ=�o��������.�p���夝J��-��c��6�8T�>$<v-7w#m�T�����Hة�����,����$g�ݪ��&x~a7�FKs�����'~��S*VX��ЎD��8�\T�����U�� watl������Bg��q�lB2Y	uĤ�C$���$�!JK�ҶC��{`��k���;D�8%�qo���x��Y�8p��O�h�ٯL�� �N�	��O���d.�?Ɓ�2j"ϼ�S�p�a��/O�U�|�R�Nh�����?��zy��;7Z>mV$,�Ҷ᲍�pɥ��tZ�R��D�9���9���s�t2�@Nm'������=���y�X(z	�H��LrY���?�����z�F�O��O���Ҹ;���Kh����6pf�j������b��^����}��H�iB�_�I�t�\�of�aK/�z%��R���'v�+��$M�{�[�i����cG��V����C�e�.O>Bsd�PGF&�f�_��8[4?�<�Wm�B��>��U+	�fR�˖���C���I�T�L۱���f./,��O���0�����O ��fc�H�v-���������C����p�#:I �Xq��0����>e�)����x^�&d]s�� �ʼV�l�"2b���z>6*N8������%�9aA"�W6̝�"	LDl��u��I��Z��#��x���A[�j�+!X'T�Ĺ��#������Ci�G4�L�LK����C3�-�.�]�l�|�zѬZ��K����vX:�?8��Rz��>$|�͒Q ��4��mDh�];=�\�H�#Ɏ5E2�Ah������.��w����_�����C����s>�POc����{�::�ّ��v�ƭ�����^��pw����:u©ח5�Iv�-{��l�X�W<Bf�ʕ�[��[�j��ࡽ��w��j�g�8��&�D=i�#E;q���>=G���;<}���Ԣ�
�(��d����pO��� A{�yal-�z��&��l�'{��@��=s܋Y	Eu�W�OU����1���S�S��r˥���Xp���h9�È�j6象<���pp��.�(�' ��LZ���'��0��"��|
��tE�.��JHK�秢v�`��D5���`�����/x6�9��<6w��-A��P�L��\_���A����~e"�MO$��:�*�#~r�>ƃ���ь�������j�yrc\Փ6�1��s	��kǕv�5��j��UzZ����m��E���T�?�ō[-f#'>%! tJ�D4e5Ŝ��F�&un#󙪬R�Kb�c��.�?5��Wl��ˬ���{�.���3Y2���S,�j��g�-����;u��M�pj���!�
�̥}��d�F�%[�z�}���3�(��O����W_����w�5��d"c�C;v�U*i�>�?Z��o��J��|���J3FC����/�뿣ɲ��rQw��k�^.���3���g���&�!��N�[w�@Tҹ���Z�Z�}�����Lg"39t���+����dI�h�	GlowNt��elr�)�S� L�LS�js��M��B�@��	L������|<;N;@\8s��]Ř�;����u�������Z|8��9�g���|hͷB?�t��Vu=5�x'��8`��6

�$�D� "N���-���pή��*۱s���-���IZ��0Kϲ��V���Kl����9&��F"�0S	s�k4�.ؙk����	س~Y��]��Z�R@�,��s���y���X.��cǎ����HФ�ܡ�G����ђ}��`���V��Mh���
��8c�8NG��,��d�:�������u��/~���~��2;ܽ��Q�=��C�#v��	�V3�w|Զn��5 �^�E#'��@���h������{7'�ςB�g���� ��M�$��lh�%%�g^��z$��������X�Ƒ�nk��ˋ����
� J}�G�$�86�\��X8/��:G�XDu�0�Rܚ���<�� :�%���c<�7?
J�P��&��͇&L������A�����q��=T���/D8V��!U'+�9���ޔ��܇�D$�p9�~Rl�|#����(�-�$�Ph���z��Λ�q�;
��}�9��7�у��
�]�H��
��$jhZڇ�==n��#v��+lێ+�Ny�l5/�l�U�d���]`۶�Z�J�9�T�lg�J���|��]wOXz�e�4��p��)�֨ΊR��l�)|Sp�(}}{��o�/��ʵ.zz��Z�!�����Xɞ}%`����Y���5��5�N��v������T�`����f.�3|�!��-g����ys�X�������֯_i�cC6<�OF�����;f����l�n~ÿuPB�S
�pO@�C��P,V��͌_Gi�L.jD.���E��M�qPKT���'�H�~k�S�d�3}]�E�I�[O7���9�����Y��<_��W-�kw�zʣi�_�-Y��n�G&Q|7��MC���p���h'~2n}��@��]�M!�F�6 ,�	�Bgr�+�J4WsC.�6s#*Fs�d(9�$�(d��z:j���J��C�b�K����8yk���߻��.�8ʹ�����.�}>@��%��`�'�7�}��1��_�mۖKm�+<�'A�;B=3yk��l�P�9�ث^�+)~����~b�� ��wMT��C2( ��)�>�$��K��`�}�"a�(
��=��7��3ms�̲��38m��y���#�ldt��O���ڛ�g^{�7�yv�>/��E,+�e�o�
�U�L��J���M7��n���f��k�#�$h�,K�?[�9WΟ�S�m���������S>�Z`�q�UE8A�
y9���'��aѱ8�j[��U+E�7��P�8bV/Fez)��ى���s�mx��>�锭\�ܖ-_9�����_�� ��r�~�~�ߏŷ|�R���W��Lԯ��"�І� �z~�w~�#��}����&���f�`m�	�6�h� +?Q>h�,|��\���&��1/8e��XlR����1�jnx6Υ.��k hb|$4$,ࢱ��D��I��d��q�a����PH�Ї�}�O�����w�r5xq+%Vx?�k��1�k�߈�Q<7�w�>����V�h�t�๰4�o���PP�;���M�>�a�C�#Ը?����Z
��x�� ʵ'�L�v���lTҙz�����_��.�b�7=�륚�sY+��R���ZmX�FV��Q �RX8��t
�>N�5���N�@7���ظ+����cL3醝���s'm��Y�JH������1��=f#�{ǯ���`����}��}Oa�Lc�-X��/���|�L��9u'�F�J�Zd��Kv���/���6����s��SO��J�FTK"E�� �,�]���;V�dTT���Z�1�p���lf���" �=�7��b8�y�RqI�L1���U\@5j�*{�?B�\%3��,w����96^"d�b��|��X��
�޴���}b�R�ģ~�	���t�Zf��t����h��i�X�� �u����ȣ�� (m@J��!c��� 8����В�3�X���&��y�&>;Pо8_t�TH�iL��9<#�}�K_�,����0f�a9`��� �`��B@vZ.�l��=�Ԧ�	�L	`ʈ`Ma8��J�v��: J�φ�2�D�!�yg������.X���˚�3�Y�Șk��z�|x�3���5��FR��Nh#��yg�@�E��q
�yE��T�a�^��d����d�$�����V�|J2ac�g-�M[��4��z"��(K��-�J�*�/{�$<q��dv��T����xG�Sy:�8S�R�(41�˹0d�iPT��[W{�|�z���(�uKeӖMe�\%���i۸y��[{�c4�_�K�7���Tz��;s�����}ph�]2��xs��HZ%n�<>:�����z{���R������������������a�V��׾�&K��zł����U'���bƹ�4���'N�t�s�� :6��<�q�8M��mu�?q܎�v�?�%��:��L��600l�t���B�
��X��J��:c+�'��;�t$!pQ�����fuL4� \٬$_1ԭ��"d�D��%2�1@�ط�9S(>*��;0�h4"���k<_���ƕ1Ҹ�a��3��x�d��0[��b�)�E�C��*j&`I�c�I`�d/4Hx`@��[h�p�1T�7���������h��8����XB����.�hu�s�?����ܯ",5y8�G��p-|Mh�{� `�����u m�lƁ�&8l� jd4Z�\�5�����>��D�0F��%P憹b-  ����IP������V}��k�9s;�R������V'E��t�=�6o�f�k�v�Xs)��	�60?�G>�)�(�x�b����%HY袁yO�x�޵Ò����{�g�'�ǎۙsg<�c��Ev٥���l��n��Dʾ�������}��E=^�IF`:����|AΛ=+���|s]w�5�������>�4�����uk-QoX�3~�644�?4�o��f��h�y�r�ı���h"^����ب��	��ھ瞴3T�L�,��Y�R�Q���t��C'�������^��s�-[���5#��Bm������,b�n"�`D''�l��e3�b����Ip��Izcs#h ����3O=�&36r��9��	P#�µxv	�x������2��46-V
�E�/Z4��D�V�GQ�G�]�[�/�����y��Ra�� �x���&ƀ����# T�z�k@��X^��>�4��LX_<'�������1h����'?� @#��C�@� �8�Ʉv��������Zg�c�Ag�8?� gm�[�_��`�P��(@�o|��'�SZE�fj����P��>�4���2|�N�@��֟���x��/Xb7��j#i��:���eg|[<t&���½h�B�19�qd3��#ㄦ��\'�(w�wݾu��!��(<pp�����  W�Zg�]�622f�]�큇h��W~�H�L�3��۪�{�0�h"Ж	�$������WU�^6��ѱ1���v���kAl��,Jܒ��F�q|��؀���������`)@�xDJKͿb��>j���d��5~*�B��l��=���=aC�t����YV����ޭ48����Dҙ��>���'lvx�
`ġ���O�k_�:s���׿�5��W^���F������.n���ccqc(�l,
�b�� ���>�FT�]���VZ/�B�)�/�e�h]���Q��SҘ�8t?~z</c�,nE��,<?�����C <�ll| Dƒ{2�h��?����k ё�aJ��̀P�3�!<?���&c�u��6�;� J����F9��`y�����8Xdj􂠅��:P�Xm����{� ?]�L������"�Zh���t_j_U��^����Y&I^J�Ն%3Y�d�FƊ6{�|���<0�.x(:XfШ�?�K��p_�v�ڭ�[@�yG��S�>���������׽��8j���A��j7�(a�"s�\�H��������w��Q$*�MHw�O��(�\🦍#`Ƅ���h���h�L�Wl�-���Ƥ�_D�@E� �*�M���j`�"�p�hЄ=)a���Xm~�v��ΗҎqJڧbGz���'���4�Q�!w�&��p�){��O��%�;�Z��V�p�GV�T�?�@ |�cI{g��n�J���=������G�,Z;|�-������Zԓ�?1�)��q��c P�u@T%m�t�����"���wm8�ņ��A�0�r��@��.aYO�<��q�D�@�BQ>ʁ�'�O�K�s \z�AK���|���s�m���#��oG��G�=���Z�ǃ����f�l�a��5�X�PwX�� �h���g�0( �\���u�څ�йV�� �=��P�Ϛ�jb,v��I�'��xX>Z��͍����f��;��{�r٤U��z�z۱k�%�eW�Ru =m�ɜG�\�y�ժIKeڼZ�C����G���}��_�E��G>2��b|�g,w���*ժ��,T栽c�]q�+�b^�v��x��G�`V�Ç{���r
S��N�
��gl��t�>��,2@�	Ne��F�*e�1Z8v���j�}#��бǩK��Y���9j "�z�$XR��?Q�BB%�[q����lxp�FGO���i�}(E��s�Ġ}�[߷ᡒ�ۢ"j ��UK]�F�i��cݐ�Ef#-���/~8e�Xo_�or4B4M VM�т�� 6���骫� �	�-	m<�m��;(��h�|�8��8��^e���f���]������N�7�6�W%P��`g�a�+GA�E�T\�(#9|�;�׀��g�~�%�)*��b�������}��|:
c	��Ppli<*�O
��u�������r����sq_���ZQ�@�J���zrT+(��eMqM��g�r��8^TG���O��Zͽ~j>� ��)3|[��v�����
۱sS��e\#�?a]]�mΜ%��5�/Yn�z����?�L�ӗ+��>�G���E@~�w����)J C�bY����)6R��1    IDAT�gfnU�;��f�%B�#b�����K/qg��X��A7��SKD��{ǭWy&/:���?s���;��/Ȓ����'���ظ�e�У�^�s/��p
K)Ւ4���b6�������ܤ~�m��T��tf!Q�`J�oDF_[&�)�=m�O1_'���#>n?�d��H[�T�K.Ygk�E叧4�X�{ m���F�n�3.�0��~�X�[Ex�A�Y�߷ϳzh9,l�� F@���G����E�1D}��|������A�I!P,a�Q	�ph> j�N,5Ȁ�����>����.�ڝ|xfq���tM����a�����W�ʩ-��+?s� exVh�2��zr����"����uO�����&|P�z��»�""�k=N����h}��� <�ƃ}��%�����; ��<�s4��/^Ѥ���h���)+m˖vݵ���;!��x�ƆKw��+�^��;��A���{�tųR܍����r�{��`3� (���r�χ��KOF9@h��e�q~'�8B���3I�����"��C��7�֚d�f.��t�Ʋ4�x�ġ�?��g�b�4C���D9hCiSPd�@5@6/+��s�펅%z�Ο�:U��H#JZ:��.^�D���{��g��+Ke�Xo�I{��ld���Od@�l�b��}����X;:�"!��c����B��[�0�<!nJ�
5}Ox�{Ȇ�����������T�V�-����t�{7PÇ�P����59_�V������\�MO�)`h*��s��
 6�j&XQE����_�U6�m��6��::8Xq,����/��}�����d��<q�>��(×���d�9j�� )�IYq�d�/��V��l�R�uJ_e����q�6I�����]�=Y3�j$0���Q9q4�tsnTc���3��?O��1g�k�{p��-{n�����`���y�����y�'6������U(  ������
����� ��V��  	N��h��4�G�U[.e4j:v�:�Uk�3���}���>j#cD-D%�q��\N8be��Sq����.���=����*m�����݉R�g����N��V�2^i���xL N�WtL�M�gCX�D_ hy �)�ĵp�J���j� /Z8<59��f���¢t\_�S?��'���%�-����Z 2
��jG7�waX_3�s���]iU
�ў1�
��ϛ����q�Į�f�%K%jV+���ˮ���7Z�Ay��[���(�V�|�#8{�O�O�uwT�5��=���DAE&)���Y?-�gk#0�YPJG���r|�N���Kj���{�ǳ��<ON硝�x ��O@��������ln�"�Z/덨�U˦y��uz�z�z/�l�͝�ǎ���<�Hk��zfŲ�����2�3n�ieq�}�t ��C/8��Ǌ��Xw�j���CZd�I���55�ԊQ��6���e��qܪ�W�O4x��AX�i�xm��F���vQ/� @j
�ć�Q�ZΓ6�spO��p�S��X�PS�<�P�#P>|G�?�1 b�1;��$!p��_�z�mW����N^���-���s�c�ev�u[�V-X�Q�J�jK���U�l����6^�z���N�d���8%ӨW�?������#���M�ɨ��9�J� �&-�����?�9�?���5��[&�:U&B0���⣨Y�1��)Z�`�B ��p���BH��o� ַ`c#gll쌝�?aC�#�6�JS5Ǝ�L�?U>�5����eQ�H�M��3�ȑXuax6��lt>ߩ&>�X��H�
Xm(ƀ(�ƈ�_Xn��f;P��G2!�d��A�uE����	��P�#A��ɠ%f��!�SA7q圏��kh�xo板au����;B��@Ӈ7��z��Kr�	Łkആ�x1�J?�B����ի�z�o������`==�Q���]��J۹�
�L:a�j�R�v[��޽Q�\M�jn@����I�әk8�H�'��"��d�b��6�<Z&�|�=�|�%��.�{wk�֙��/!p���:�VB<�ł���'��3)� 4�?_�����R? ��؉���@�Ɔ���G%_R�6;�7`߾��Z�����4�˗��ZםJ��Z �@,*%0�|h�Ӂ/K5R�m�iu>����ب	�H�Nw�l��ę�6���G�����P���gW�>�V�6�=t�J���S��r�</s�ld���Y x�Y�sg<%��.�v�۸/V � �Q��t��O"�_ Z����45p��9y��7�|��X#�s�e�u˥V��{�b�����*ik��U=���*��oo��J������׵�����r�7�H)�\���i�_�������6p���!�4���F�hB#�nr�'�جh�a�n����q��4K�-�"Sr��������8j�Ҙe3˥��]�;�w̱#����S�BUh�+����ΪY��C3BP >��je��8N�p I9V�ĮPs
AZ!��C�C�V��i��DA���y���ID*a ���E�*�F��(,������~;��k����s���������_/�!�}Ё!�F�^����?����ʃ�k�`~�����\��������f��A۵�J���͖JT�FD1�n�u��x�f͚g�]�j-�-��p��{�R�'��:�%I����)�p�7��LE�|&���[S>��(��S8|��帝��A�C�h�>��Xlbi~�z�@��V��^{Ķ��mլK�g��Jy������j%��LZ[{��}��~�)�4)V�I�'��B�Oʣ�������y~�a�TdC�Zn�y*�G �	7�+Q�l�i$����xEIp�q�M�Lo�O<t�4q<����&��$_ׄz�2�Г%#�E� �*�;��է`)�@�yF`p}��*Ĕ��0���r��B	��@l���.8|U�'������s4pﵜ[ӣ��o߶��ch�J8��Ixe�f�����M�Z�Y"�v�8U]��'�G=�{/�]ȘJ�z��T�P$T@��iGd����i�}��}�����00��(�	���&�\0	/c�jz�5e9��kG��d�h��h:m��wl�*�#F��$��g�R6{����B��J�l6��˩'ν0�������J�*��c�㈆�����w�C�1/p��7p� z�(+��8���y*#	���&�Fq�Y(Jl��⚊D�#Y��r$��g�A&6�|���0�H���r�9��W9�0�D������h��=�x��(r-j���h�{?�E�,���Y���,�oV+Y�2�Y�:,��rw��/V�\JX���L�ݪ��er9+�"���~~0j����z�S����d�˼`�[����jg4�O�O&_��f����K��f�vv���8<<��ZWW�'Zș'`�����W�� /i��AܫUy?-{��{�"�4j$$%��5��.�'��L�#3e�j�8Y%���w`���ݿO����
��^@4�v���4v� E,)��r%1�/JbGCb���K���`��wfgg��������~��eؙ!�/��s]{�Ιs��y��������4�dh:wx��܇���K��s��P����9�D���}�)��H֬\�bi�RP�UK��̯Y5V���M-�m��,;P�Z,i�x�^ۇ�<�\32���*cS�L���W��/t"4`��ɣ:�.0���
:=��9��������Z���}F��?�����2|�s %-%_{{���'�oނ��h�bkjn�b�`'QX�����>셖��Z��mJ#`�ʙ��D��~�]1�p�Q����G���?������Xv���ɘ�ke��b:�����%;|�۲y4#:=Ǽ�ϼ���/����E�PE�g}�$�h<<H A�?yF�=z���q��#f���>5/�]�	�36y�Xˤ(�V��Y�,f�B��?�.��f�B3���h���O����G��?~ꖺ�&�!�o~�o��@���������&3]rT���j����cC����Δ�o�׎>f�==~��Jf7π�?|.�?yʤ�x�?=t���f.$q�������
d�-[�£+H�bQ�z�=�ڹB*�&�v��qkۿ����7<2m=��"�H�!,��pp�*� �?8OTI�7}�fC^��}ʶkףv�s���ojL8�{נXʒ�&۹����v;q�ߒ�Fw`�@�3;������q��#N'���E��f�Q:�
N�@[I8�
���
�g���
�7=Ŀ�ᛈ�l����v�RkH�;|I��KY�T�ɓf؆�[��D�56��8�b��e�X���S��)E��:F�i��!AHTAx.o)�''>�/k�3?c�L��!������d>�
�B�f��zh�}��o�B`�ވ����G+�f͂������R{�e/{��$9�6V�y�R�d���8���9,�xZ���X��O</U��%�0d�ǆ�4.��i�z���ݹ���>dU��J��V��KZ:�b:���������[��٩�ٳ��O{J	�����U�S��M�ld���#����B��X�N��u��7aȹ�>Gg�4���RD���5�ym3���c�u�e&��S}�y�_d�
��)��i�4y��=4��t`8�u���J,@��<���=���(�¿r��J����`-#jzz�F���������>�;u*�&�yt�����G+�K:"Mq�^��^��ߴ�&
d嬘�z�*Ijjij�~!�7�_o�c�Y�q�;R�i��z7����&Fm_lJ�aB�9��C� 0�}�$�{��>��������:h��)��oHc�P,Y:�jm{=%ɋ����-��>8|�?R�/B���Ĵ��8�t�OC�ۢQ;Q�����}��Ϲa�7��S��$��F��ty���+�T�ui��5�wcV,e��u�57�؊U�,f��Oo(�G�m�稱��~��?��p�(@�ƴ'e����Om��Paޣ���D}g���%���T �����jժ-\�ȦO�i�M�J7xe�}m쓟�����Y�q�uV�>[�m�����Z�
�8aV������������y;�^{��?��J�R�FsC�]�b��^w����$�P7 T�=��s#D�j�rS㇘a�ˡ����|caRu2Z�-/|ڱJѱ���tٱcv�H��v����Z,D, ��=�e��+���T���s��
#�w`c)5D/����y�_�.~_a�}E��2Z��#�����xN��������>/�y�J+��M'�&mN-=�V��d�w�
eknj�dH�:d�!�1V���GA��د��Z��l��	����G��?�yg�r-��|[6��B~����:w����}���㌍�0�^��ټ�����Ŋ��=�ȣv��
�CB��.�?i��t�m�������xOo�ug��B�Rɸ���/�+.����Az觶{ד�L%,�ΈU���ռ�ґ�ݶh�{�^7�%J�I��ۭ�B곐�T�;������g�d|l��r�$��/@����U*v��k߷ݣH�u���{��6�CcOz�r���>Ϥ��(6>�����ƣ�Ȅ	�|N��Tq���F>/:8j	����C���b�97�g��v��\�_m�<`kW�g7���d�j�l��O�j�nt��n2��3C"��D@!��By�������
�l�r[�q��� ��@�6
UpaB&|���|�j�(��jκ�qő���sߙ�6;r䘭]���ѓ���n��K_��=��9�i_^�u���oV	�ل���}�-[z��
v�}w۬����T�:�a�R�q�%�iJ��;U�W��k��/>��� �$qू#� :,�Ph����8�}Ī)K�O5k�N򪞅b�'�466[[�A�����=A��@�ޣ�����o�z��$y1.�K'�W��;�E4u��te��2�yM�bcC�\�9{�e����h��%���=6X�9�ۜ�X��6oZm�*��kV+Vm��%6k�*+V�V.��Z����ӂ�G�� ���G�b�[�ƌku*�� �3�u!���T�_�?e?8�rΎ����`:;;,I+�xh��Y=|����g-�/����fϙg�x���;�5(���>g��m��zz�����[�O�<���G�q���������9z��zp����w[��#�y$kK��R��Z��7�<�4C�P��B��ҡ�����]��<l$6E�p��覧�l�z��b�͚�v�H������}��W,a�;�����S{��X���i��U��x�Ё�+_��]r�e~ppӺ񢋶�&�l���/�9�a��&�.=CY�r����-�0�c�S���+���˸�r.��Z~*�B�V�a-���/�t4F[y
��U����������*�Aa���>����4�Ud-���I�ɀ��i�pMeG�*(�.c>�x����E!ߌ�M~�9�����-ާ�E)K����՞Pb��
���p�O/���f�b۲e�U�}�L&,^1�>k��Y��*��b���:=s= ��Y苡�B�����2&���y[�]�W�������N$��O'?U��_�����'��&Nh�	�Z��=���Y�6Y6W��;;�RK�ɓ��v����rNM�O�3�x�VXt�G��,�}F�PՒE�?w�]�u���>�����]v�k=R���C����fX2��S������i��q�V������R�'�:��fs���OO������'�����r Y�7kH&,��Y�������;݁��4���uڽ�?d�\���Й����z���ꆍJF�a���osС�O6��m��^@G/V�OMz� ��9P��<(<T�) ��-0侀���h"m|���(�34�@ 
K5v�q+��ļh��V�ͅP�ƨ�`	�A�Q�ƭ�b͇~�<J H��Ґ?�s0^�c� ��:�� ��
�1N֌9�s\�N��t�%��4]���ֽ���u��C���D��*�%�,0"�O�흼���7sQ'���%��X��+ϳ͛WY��o���e?a��]��;y�����/��͵r������~��)g��⋼�<?
g�fCP��৒��g����}������ov�sm⤱�c�ϭR����l�v�9`k�����\���B�x�����=%S=j���Y���>���[���v��U��@�}�߰�/�`�X�����p���Y;r�U*��v�5L96:�ޮ�_�MMo>� @�����}׭��8��u UR*��%gt��J�����}����SGͪ��h0��X۳'8|��g.�����!�s�h(��h'����c��<c�={���;<�B~�֕$�ѺR�BQmz(�I��(xHs�ʀ��F#�� �� �!��Um 	"��Lt�+�O���{�nc0	��J{H *������q�"� �p��B�u��2~=�,�cM�^�F[����?�HT�%��c�\SV��������e�N8��p���u����+��P�!��6�X�p����o�8�4i>��x�ɚ�L�ISfz#u2���N�C��g7̅yt������-1�G��G�O�'���g�+�K�X��ڳ�q{��o�ʕ�l��V۽g��$��Rͪ��=���4���'\���
�U�yٮ={�'����G2Z��Po1X�{�����?�^�ɪ��>�����L}���'��[.�#]�A�G��ѡ��,"�J
�PP��8|��l43q�j���<b�o�`:~f�OX�T�LC4�x���i��費�}����&�T 5�3O�����P�\�4s���6���^�!�P9\�k�6����0c#���)o,�|G7�6�4h��@F�q�'j�*�,��QPR䖛�ޗ9lE*�vQ�d���
n����S��PU�b�    IDAT ƳH;}$@�΅��h.���q�
�|J�������o�;���X��yn�8lֆ=�ƪ����T9������2�%$������{�{G�uGC�����z�۴q��q$��|�X"�%�s��G�<�"�z�,I"g-D��kh��]]��=�Wu@��8;�[@YC�!H�f��e��٥p=����<��~������ĉ���m��KE�R��lޏ��w���2������A�����mFֽ��9��w�?�GkK����&O��η�n�S��Nul��D���T�:1`��d��/��^�җ:xP����o���'u����$�:����k�7��m�ڑ��<h����&;S��//��'�#��,�Y*�|$�D�G�9��I^ݧr�L�X�Z���9�3�|��_���_��_ٛ��&[�|���b��Ǒ��9��	~e/+�M�T4ę�( �
�J���h��p@�4K��z��4z(��c�gS�(W/*Jܺ@?��.!%zHt��*����BF 
�3o�>�����{�y�% ��2�����.�2�c�ŵ٫p�\KN%D͝Nn,��O ���Y@Q?E�ϴF<�z\h=�N�g��O�{�f�qo�N��WY<^�r)��=e�c��/k�c&��/~��*���O�;�D�P�+����i*���Y"�A��F�'��g��|,<�����8��}�~t�]6}�8ki�XGg�ˑ�PW(�~�C��ȱS���o/x���+�\j'Or���/|�N��v��|�V�YL�����&�P�xʶn��^|٥��sº�:�����8y�ʕ�%q+{S���c);~�{���&�_��5N�pҹ��ˁ���~���XhWl2{��A�_u���=Z��r6ƦM�BM��7<C$y��8j�	�$k�JIgw8�c�δ؎���;��;g�t�K��S�'1�#w�Ղ�O�UW]��� @���w���C{��"��j���E]��1����-��0�QJCܺ�n6���Ґ��^`!MYZ��q�9�w�;E��q�v���ʚ�`":F<u��$Ǯ��k���`�~Y%|�W�bQ;r���FAC�X��`3$��0c�,9��ή]�|��@�{I(���[ȱ�Ϩ7��G�,YC�LtMt]~
�7/��:�|:"��×f.O�}��_��Ų���CSC�J�|�y��Y������V/�\)ǩ�˜�7n�;~�~����zg�@߲�?�я:��<+����}h��h�����u���u�ú���l�+������	;��k:�X_o�^�����f�2v���; ��*hρ�(�݈v�I3���׿�Z�Ҿ:�ڮ�OZo�)KRʙ�o޹'i�J�j��󗬶+��!��D�s�{�8�}� ő�/��O��/��n��&w&�Y�!g�{��(�U����W�R�Y:�D2f�b�R�F+Wv�D���5wX[,f��p`f>��>h+��7�!lj����r�']�|�;��!��gy@���A�C[=r9(ꔅ	ˋM�5ѐY>��h�(�A���|>�;c D!�!�9�X�+g��|0���5U���" Y'����Su��S*Ғ�{��)J�uHj͹�"���s-�s͘��s4K5|ѳȂ���]�z���&\�R"��s��PEX���H�p]�IT����v(9o͙�>��Ng�)A��D��(E!���8�-K��J`�4E��.�8�O���~)�L��榘�C�D�O���|�i��U��(�@Ѵ�eZ\�O{�>��+���A�_��Я���(+KJ�g���I<���jլ���i���Y6G���G�Bɚ[-�/{��qc'��������;��A��3ٔf6jU�xh�H]Up��ۅm�9�j�����O~�#;��a�b�-�;ޖ/_a��l�Y�X_߀o��[�V�?8|�q�I����?���]w���x<l��f�\(���G�;�k���Y���T�fU��d��h?GtO�,��д"�$V%���U=�|F�d<�&Z?4����N>�ʳ~�S��tTϏ��\2� �Ќ �K@�"��B`��}��ph�'�y8�&�$� ,�.-|$��0�9��LBp��"hq���c�)��cf��G)cz��\�3�G �<��3���Ҁ&���V}���K^����p/��K#`"K.v�ʘ��ʕ+]��pD������sM9b�����d���5t$��{�;�\��9���5`mn|�y�����x������e�l�B���`�����݊�8|�	��˖0�Eђ���b�X�
Ţ+J�Z�&O�i˖��J~?�%�I���Wc#M[ʮ����u@�'�����W5n	tYV�=B��[�E��ﲥK���wn�n��~;~�;�)�BH�̙sl�ʵ^h2F��Z��o_��/��t��s��!0Z=6�Lu~�u��i�F����Bo�́�����k�X�&L�ds��3/�M$~,�& ��X���ȍh�lG�I�r/�o��o�q*�tp�}v=�����I�Y�R�)B��ԩ�=��V��_f��˂�l��V.#��8��WB	�fӽ�5�sڈ��9�����;�0ǯ�إ_��W�Y8�D(���@���>g�|�+�
 ӵk�:� ��CMH�A�O^UNB�+�xrσ%G����kD�5k�g��0gPvX)j�~�m�����6w��hx$��A�%�C�@C� \\��B����"��p=���q}� ��? ��e O(@+ׄ˿���z���گ9@�RB��<@�#��Bp���[n���F�+���A(�,W, ��A,� ��]����g��,��3��E���������}rMX#� ���`��=4[��ૈ�D�)�oO�2|G���[8o�-]�Ъ%:��=I���R�f3gͷ+.�;W�����)錒�X����=uʱ��y�E���u���/�gy�����\�
�8C	y�k_m��u��\(�Ѯ�v�P�𠱡�.\lc�O򂊍MM��?�/�v�ϕ�h�轢��^�4����$+��~P.��W��!�6��M�ߟ�����������?~Jq�lT6?}aqS1�
�\���_�ʠ�)� ��X`��\|z���_�O<hǺ�[KC�J���ͦ�Ix�۾}�=��G<f�B�C�jη���
����C����׿Ձ�g��׾fO<�sOhan���@q��!����t8�� _��v��)�2�4y@Q��p,�\��ܓ���'�=�y�s� ��.�`ܙ�\�w�֭x �	5B��9����T�y��b�/�uh0ƈ?��lXH 4���S L�}XX '�A���l�F�'���	��!8s�<#τpŢ �����ٯP��9����y�#�*G�o��o�}X։�@�s/�k�6�����,����1�&�N�}Ü�̿���ꂛy欈Fb��'�)����f�G��h��v4���Ϫ��m�ƕN��I_��j�wĬ�e��]�Ɋ%B&���|ɝ��7�C�;��n�[��H�?a�$Wz��ST${�3L�?���Žy�W��J�9a�Xߋ�Jy��Q(S��[=���;��g�5g=��h�6W������ji��0O��!�K���D�������^�>��x*�>��'o;w��~��v����2�i�p�ho�xh��o��MZ �D����}?�
��hh�̑���l���Б���Ү%KŃ�_���j���{~�����=�B E����B��ac��‿�s����::� P|ի^b�=�<�����h� 0g^8$r2����a����G ˈ�Vh�h��6 
��ÆF����%�!�   <րC��"Дo�sO�t@��v�o4~�eВ0P0��� P�V��r`�,��5f�h�h̀>ό���	B >�3�@�4N��5��'�)$F� ��AX"�����Cb1�>�����D�p},&����A�#�{"`���9�^��.�'����#9��� b�y&4c��Dp` h�OΎ"�$ ���;|)�P,���5K<cߪy���Z�a'�P�z���u[,�i�r��u'�' ����?�1����,�ٳ�z�7�6���|�c�R�ϣ\$@�yϿ�.ܼ��iTidM�p��v%�$Mŭ�ʺ�w&!pVW��b�����y�p�O��Or>�is�Nu�9cƌ�C���lX���~Sf�Y��ϡ��&����CE���� ���Pa��4��p�n�R�֒9oP�]���x� �}8�2��,^|�M�>���G��PB[�N���k|�2'X��O��2�(���������{ #a��|̫,$@����3�I��������Ƽ1���
���so��f
�:tȅ��ڱ�rJs]@���1���9�p#���c�q�C�kG���P"$������=� �'����~ m��S��Oh�B����F�h�PiD�(D���[).�`yp=��8q�<��ڡ�h�X8�)��E�@��B8 �/��s!�z���j��=Þ�o�`�Z@X#@x&�-
7)oӦΪG��9ڇ�ΔQ�$����R�Z��W5|l)��B��1c'�KVX2�h��R�Wt���op���|��.(YC����}���d�27��!�."���f���`��R����B��X����ΰ�E���Z<a}�Hk�^g5�_~�����j8�?�$�v�"M<�B!;�~����t�oEˤ��TZ��B��_��_��Dy��C��h�����-�q"z-�x����U=���Wky+�؞}O؉c�,ӀI�������j�,�ޤ�+$y-�3��V��h�?�q�$y�I�1 �}�� D��PCc( Q�Y/Om����������I����Y��]�Ce�2��e�?�C�p� �	x�
#�@c:s���4n@P�|O��1&��[�L�#��z ���@`��h��A	N\�ﲏ?ό Ch�>��2V���%��7�G��X�D�H��3
I�E� <PMF@]{T,4�dyvE�)Z�9�|ȷ�ȗ(��'�s�gB�����{�L�nY����O�����5��zl��e�y�*���Z�jD�4�،����ɳ����C����k�t���y�5��S�7��>*���<ɡ�{�_�A� �a>�'='ק�K�ۛ���!D���+,s�9E���r�����2���=|�]񩞞�7�nB����Oo4B:}����K[?8�нG���f�)'���q���9�8���X@1���5�{���G�R�Ǣ����s���ai	�fh��n��v��S������>ف��b�:�/�&R	����11^LN�����(h�������"��?h/4>Q��h��1�����%=��b�a��
	�o
)0E�ֈ��'�(��Xt��U�d�H�(�C�T+�� `|Ou\��>�Z��\GQR$����r=��M֤"�؛\K�+t�g��*���r�!���e�!D���h�|NJ��#d���?`�gEI��<p-��n���:��b%p�}��i����y����}�+�АIX!�m�/�u�.���_�ڤI��${*=�jP<��;�G��@�<ɋ�?
������8�U	���U���B��u���@���38���8��h>���i���@Q��4�)�&_{��f�������I�����fU̓<�0s��җP1����7eZ���wP�OA�
�xk4A8Mi8�������>��G>2�@h���*�v&��"a)KZ���L�b]'xI�b)�<���?l���'^�ڧR�;(�R��p�����p�vc����b>p�AO *  �Qx
��ϡBbJ����7�����[U�l\��aN�	3~Ɔ���@B���u|�4~w��+|
��;��X�@��*?@Bٰ��W������)M�����ݮ��{K8z_龾A_��q�����T��br�	�
G2t����N��!����G�Gs%��s�̫���{�4����SF5SM!Q�Q�$���[��8^`k�,�t�jTM�C���KmּU��W���d2�)-$t��hL{G0��sS��O����� e_�w�5�Y��`-�|� <j�� �J�=���u���zC�
�J���B)���z�s��f��m�>�����3j�5����^���
~BX.FA������]*�tS�8yN�IT�d� Lp�*(Հ���o�;~0U����UճZ���=Cq7�>5J0c2;z�ö?��� ��2����{?[�D�����/tǫk6�vc�\�y�X4�F�I|���s�� � Z<�,��CX��@ �
�s/zB�%��i�:P�'�4DJ�LS~���e�&d�E�1i_|A��4Ƭ���"��rUn�������wyN�/��Z�l��D�B��A�/E���" x�Q8���e �������J���a˜��+!-Ag���|f(x�<����tV��Z�B�������B��p���S$'g�-�իϳT�j�R�
��-\����_c�J�2���C�Fē�z��Ԩr>��W/G(Z=��,Z��!�'�H�#��u��ϧS��T=��s���)�����M'�<�s��030�'b�$n�
�w+�/�ԁ{+�U�6�{��O&��4�W��{�ő&�CqzA��E��u���ٗJƬ�����s�>q�k�P��H���G��w�o�Y��]F�9#��� �5�����s�n��R������C��� �04�Q���H?��<#��sv�P:�kp �� ��f�=_A��m�T���z)dt@��ӜųhW�\h[6�6����)U-�j�9�۬��󗢇�r���p,|����`�̠q�T�,�`�?���*��n��di5fBR�W�> i�I�=�B��C�����ʭ����y�p��B�	� n�bg����!rE�* ;!��<�B�������H&��c6 �?�hrI��a^����:���O�c�d/�J��il����=���
�PŇ����_d�f�䅹;r���ND�?��NJ]*�ϸ���,����m �_ڰ��у�\�g�5��'����/�n~6?�pc{��O�R��{�nظ�jeJ9Sч�кcl�����:ަL�a��YS�8/�\Ĳ��W�lx@������9T`�4{�9�S�Ƈ�#�NTD�<gIB9��"r�T>���Z
V�5����OX�<��?i�|��>;t.��s���?^�`�U}�tTN�`~�<��S�.y%P��K�e�e�G�;�F�Y��l�-( 'Ǐ�P�UG�v�P���u�I��Q�J՚[&؞������C=�	Vb68�PO|u�p$�!$��5�\��Q矿���0�I�����""H�h��Eل����^��p�b=Ȁ;�q�z4ƿ����* I^O�����C3�zd�mӆl�����ސ�X�HDƊ嘍i�`7]h�<�C��*UK%3�h@��$�|��A�od�K(��ɏ�)�Q���N)5�y�B('Ih!h!j$�ǕM|�жi�Џ�7p?K�$��J<���3A�NXA�w��\� ��0�j$�}���$�37�k#̐�I��Åz�����G�\���7�-V/�[�O�l��'��{�%�S�&.�g͘�tV�p�����f�����t�+��ꡉ8��w��ͳ@-��I�l���<�8;�� 9N�{�����ϥy*�?��C �vklHY6�m�V/���ά��(
"� �X��Ŋ�3Ѷ\x���!L
�'I^|	�-�s�\�5��;���9O�����ij�e��+��R*{���	-G4}�ߛ0�&�:�O�2�/����{�i��D�T��o�+�����'/� ~P���N�B�#a!� J�@��G�'`K4�����B�CT$o�    IDAT=��5f8��'Z�����UK���֫Ikk?b?r��z�I�}p�͟;��1�	�EG�F���ybŊP'��@<8B�������AU/�+��{.��sm��טkY�RZ��ϵg��2���O=,r����CU�T�,ޒ-^0Ӗ-_d��P�Y2��`
��?�2��l����b��/& V ���_��C�dE��E�I�Q��a��b�!(T%����G
������������ng�O=���n���:���$/xp�RK�)�Q��G�"qy)|���(� Z@��(���Ђ밍�Y)"M�Q/�ŦË�
��[�Zo�I/�L�(�&V�ZKZS�D��/x�z�@%[�p�͟7+d�B�h�K8y\�<�-�08^�|@�':ģ�Ik
��B�P�gb=���2fEJ�Sʌ�tT���2��8Nk�Q�9���:���Z�2��%S+�<d���P���Lc�%S���<�*U��:�� �zb� /�y��Y⥈,�a���5�.U��AqW����x(9%"���g���K0傥����O�4����G+�P����h�l�F��S�jH���-t�pnii�E�e��,�;�vR�66��uF�5��Q�o�j�x�I]���v's��}m�����>K��?Md���d�}y�1�'��Λ�%��//�k8�G\����o
܉���\����X1��p4ro����}�=���ϊ��"�c~Jy��U3�O�����>��t�Ϥ�V*g��9f-�)�2�+18�A��ĩ�f�z���cA�S�z
0τ�=�aťpVi�Hi��E�D�Jm(d�L��ǒ��CkS��\�ԦN�l���>Ι��<�4�87	���{��4N�R���U���b��v���`��fO�m��_�9�f�E���MJ��kRH������?�I�#�H�����iq��+��n�,�pm�6Q��?b��<i�l�e�^�ө�QJ�'v�c]����gΜn��~�3F�	��|.�WQp�����_q�K9���@��p��B�3�����g����w�OQi���?3�s>���:E�-=��Z���� �C5Oj����9k�]z鋽�o2I&P�p���!ڇr�p�(e仼���p�3�T�q�?����G��	�$'f��6�lkl�0���X�ʢ{���?�'�[���B�D����Io9+9��K:WC&/N�J(�If���+^�r�0n�s}D��S�N��\2�0Ƕo��}l	o��%�dh�
� ~�EI�UGvM�̹t���JV�^��b%۽�!��M�Ȃ��|�7N�f�ut���&%~��U��G (!e$�׭e�~&?E�Q|%J��Z��
@8ʔU���� ��Q2���
�hR
�>�@�E���~r�X�6�(��CNa�<��!�\���F����I�o9�d��}�C�+�\t"�a���C��d9�"HX#Y����"K�<������h�g.f�]�|*��퓴B�7�wX�ܬ��n+W,��X-�h�bŒ���[(a!�����;`�&ݟu���6Dӕ�^���W؟�ٟ�Y�B�zq~ɘ�ҭjT)L�(��m��\��Ək�=��'�0c%8�����;�)���`��fa+4t����Z����ꎢX�3M~�_do|�묥�1X�>|�v<��u>hM�F�=w��w��:e�KUK�3��J-6
�!P�v=un���S%�M�g�?��O�#�xp�>��{��ah_�x�v�z�N�8`�B֒�%c���IKc�x۳��{߃6�������i>2����hN!*~�vv�u�ɆV�3�B��E	I@ոK��(� �����åB����G�5%PD��k1&e�J�]	/�[��響�
�IX*ƛ��B�{�:�k�\OUe��7����s�R��e)Ei���sܛ�Y��ҳ�7����SB����5�	�_O��~�O��P�t*f�B�mް��o\a�b�ҙ8ͳ<ο/�9�Z[�ٺ�<ڇ��yXl,P���Tۇ�Y{���k�[�盽�P�-@(P��o��"�٦t���Y�\�\��k����<��,��#X�����^!V�>�
�P�`}O�'M�r�Y�u�֛�{z�=S���$��y\�)S�7_�*����V-Yϩ���#?�'�|�Nv���f���/�bp�]�l��^��#` �������
�S_���ԽA�!���fΞ�%��4
�C� 7R�'����	�9u�N�<l�~zc�V�X�XC�kk;����Bm�~(��}��3X��Z�lF6;σp �pg�R߈�a�J�^�q�?'�U�+����Ł�����Ɛud>)��f�9c�GF��!sH����q]擒J����z|���N�Q�D �_�� �}d���&L|�^�ʳ�ٽ�AV�E�����B�j��{��� �oX�� sĵm|Iܟ�9撹C9�w�&*/j�L�2�+�j�x�$.�mP�_�Ϟ�<�G�����S�e�r[�a�U����$�����i6a���I�@��垓!䓤O/R*�y�k��G)�����y6�d��A������#�@Nb)3�I���K����{�b��{m����s�c�굶v�&���%�Le�;��fh���BEÿ��ugga��[?���s�3|��aH� ݛ�'o|�l����kk�i?{�^���MQ�b�jI�!�j��_�%KWٺ���9����}����)�P�p��+��~͵oqI ��<hm�G���zmr�U�=�޶ݎ>�!��$2�&ۻ�34sɖ�ݤ�ϬuW����q �ď?��mkmE����u��9�S8(<֍�u@�������=���T����>�`��6�8�i��e� ~��O:�p㾔� �ɑ@s�z����cԴᙼ�s<X`���Yփ}��!�(W�㟱"����������C�s;�^MI���O>Z!�{�Y�ʝ�	z=pO�hQJ��_��"�3.������X�p�wXc�\��&h �%�����5#y��O-�b��3|�}⵼��x�fM-m���6v�T��˚�.�֡�C2c���,}~9��\������;n�Az#�����9�;��B��#���<��`A�R�q�i{�ч��'wG�1�K���z�5���V*�l` g���?��Q3�a�
��{����m���~8�w����Z�Z�7��Ͱj�h�>���������`��KK���w>W���S��_��lŮz�[h �]9�2���� ��y�k�>��O;� ro��M�D�i�=(���?Z��Uc�I&,�(Y���־o��j%�P��\��G���)�?!��_�X-�FJ��� 	��j��@?�Y^��KD��h�<� g�	 ����e��?��?�k|��?�/�@�i:z���ŢMQ�N�� ��V��F��É��`.Y�@G.�=�3`]L�:Ʌ%�)����\��hX.T'eLX>T[���vN�̯��9�K�y���?�k����;4|@��`�ױ�G��P�Mj!!d�/h@ ����{D�QdA�r�
?t"�E��BbL������g�UF�}���)�`���Z��֭_j����9#0n��l����a�Q!��]h��D�F1���:0f�����Vk<eͭ-���WzIg�?���X��a�{�ö�\>�O2Q�#��m�欄<u�{C�|��kv���,�����~�-Xx�o��|ͅ>��|RZ�(�svk���?� �i��ٟ�ɻ��a��}��ٺ˭Z�Z[�.���]��Y���v����f�tۖ���9|�2aY�K_[�G( 	��}�{���ń�۶�,@��06�\ФG�},n�Z�j�y��v�X��k{�
���
�����q����M� -6�G4?ټ<�f6���ƾ�-Fh�@�2ln9����̛@t��j)@{�'?�@e�5Lj5�ȸ/��T��µ��i<���+!r��E�s��d��C��-娱�кyV��5�y��_�6���ͅ@���u~��<��'w� �U����b>���p=,�xz#�Rv���c��+Wz�4�{
���PE�!X<(X!������e/1G졨������ь��?���D�V.[`�6,��J/x�����Y�-o�V��{�s��sJ�y=�9m'=������s~ޒ�}��wT�,`����+�	�|��{��߶���)T�N���o,�Z��}V*Ǭ�x��ʥ/�K.y��3����ӳ�i�r���=��붭���a8��DC�9m��p���J��:q�~��o��e�������ug��R�ӝ����l����6w�b�r��g��jY|�EW�q�U���e 0���"� �5����DȌ�Ex&E���:����y�
�~�E��D������i�_����
�D�'��.~_��&��w�.PD���`i^�3���IVh�h����g�xa#<�3 >��(�CA3Ѷ��];��� ���}����چ��h� ����}$˫\)�8xa�߸?��3X*_�Hx�G�((��K_�VԞ��#�lX(T<廔�� ��Iz%�	j@����}�.όe�����)8�y߳k��=#�g>��\ ���G�T�'�Wq��zU�P�'I!�ꀭ]u��߰�҉�F#��Y���u�H4[�d0�Xܳ� tѢ�&g�g~���>Ŋ͘5ӕ��v�g�Q|��P|�s��_؋�S�'��c?�x�-_��&�c;v�E%�$䥬�7k��t���v�D����`���w{%�#�N:%�s{h�?^��?��������y��m7�`�I۷�q��[_����V.�Yǁ=�M�S����Z��C��ڎ��KVx�T �k�Q���w%�GQ��b��C�븃D����>�P�3 "pJV�����Nkk{Ҋ�^knL{)j�留�}Z_��`i��l��YV�~$�a�W\?T�ҥ��8>����^��Q�]8oh4_�X>80�<��&�"(&N��3�	���C� � f��C �e_s�N��v��2� &����ϐ�?��$3��j�O�<���������G�:S��b]� о�7_��^1����h�?/�A�#��cg~^��K��_��S��茙�&X!(<B Z뭩�ѝ��
A�傰Ta����������B�Y�*���N^T�ݸn�mش�j��OTi��V��9K��������4y5\b�CE�������hwkݣ},a�}�����7��)^�q,a�S�	5��X~"�9�(��{����a�2�8q����J�Q�L�-�-��]m^|��'g=}y����ߚ[�Y.[��|�c�Ѿo���9��O/�r�Gz�{�:��_�7
Y8���Ʒ��g���v�7���������|X�j%i}�y��+���w���e���Fʣ��������B��h� #��Vv����v���@�T��/9w��y��;rp���V��Rλ6���X�ہC��{�L�LC�
Xϛ7'���k����+�ꪩ�%����'������n�Mp�j<�g����;��w�P���] ���,%4o�V�Z"�`'�1 ,C�i�p�{�X�y��o��8��>%�X#iϬ-�`�<�Ȝ�7Y�'�{X>�=����>��<3���������+��F�0G(���w�� �N��Rr��ޔ^{I���B�OE�9R�آԠr:Ȣ B(�i�U	��8�D���c�#fӽ�?�\���(���O���[�fm�ʅ�y�*K'jV,����V($��a���0�����uʜתa�]!����٩>4�P2� ~ᅛ}MX�T�jemI�"�G�����??w�z�~t�7lŊ�6}�T{��G�Z�'/h���,�h��G���d�'n�L�����ܳg��&���ׯC���_����~�<�d��Fx������w��55��Z�ٿ��?�E�-m�W����!y���~��~�ʵ�=^��.�
�L6a]8�?��X�K.��M4/�M��p-]��7����nΣQ@���Wԑ�{T�|�������U�$%��*W�6n�4{��6��COZ_o1����m��6w������r�у��P̊� j��U恟�gW��*��h�\W	[��G��F���j��\ �\��o�D%W)�_��Z����
��}�[���9�џ�R�38e�)7@m�J@SG�~݋uT8��y�3��5ŕG�A֏��T)�?��b�?p�T��	�g!c�9�H$���O�mUP�/�BC׋�c��14���H,,�:y͝��N^�5���Ջm��%��o����:M�ן�1�&��~�R���{��J=�'a1����[�p�Z�I�я~�[�2.|?(������s*kN������g��g����1}�577Z{�^��(��T�1{�g;-�i��ǻmݺ�쥿��Ǝ�d�v����S�N�?���[g/��F�`�1aM��r�6[�v��,���ʀuu:���]����J7ہ���y脝8U�����\�����)�8����H���щ���ܻ��ݩ*f�/��hn�t���Ås�}�N�Q��s�
�>76���L|�����x؎�pb��Ϝ19�i�*pÃ?�*�#�s���f-j`E3�=Z�Rq *��<)��M���P�: #Z/��?@(�s}����=s����氢a�!�=�/�&��X
<#���+ˁ{�ys}�+��s�;�Sy�ų�󀇚�3V�����%$��3�¼���{pO�Y;w˴�V�,��ʭ���7��2��J�����ESro������i�E�:�Z�(���~	����?w�i��U<�w��́���W,؆u���-k���'E���%l�l���j�/Xn�\Ś[�?�Y�����[��Af���!jg�	��Z��BAOr�yvĬ7c���p��+���'-��B1�:�3ꊱ�-�c��?o?��Þ�՛�����S��w�|F����l@��Q�&O��K�����N�b�8�P<ekW���\s�UJ9+���c�#��Ȟ�ŇO��	ո�eK�(���.X������㧲K�����+�� �N��p��׹�@4�����pM����f6���-�g�'��b�ϓ�0)S�9�{o�=�}��lt��l���6s�3JZ�� ��p�0Y�d�8q�/���9p�lv�`����������9<�CB� �t��	��3C����4Y�(������*x2��a�������<BN<�����rc\|�5b�rƁPC�#�/������@ �(�7~|!̓'dM��kϸ���S��d�TB�H�W�>�a~� "�D@/��f�j�0�`��٫Ap�7et�������b��,C	,��>�KSԂ��W�N��ГV++Hc~
��4�o��L��^[�`�-[���P�������y���<j�B��O�����ʁ��k���k�Tj;g��r�-!(�=�S�e��Q��3�l��U�}�־�������',CK�B?��ez��6o���n�fkjn�����˭_�g��%dߟ�Uo�r����+>������8O�f�KUZj�<���T�����~��ֶw�e�h	w�,�`��۰��;���,.�@4HT{��%��F� ��c��M�1݋E�� ��!���>�i؃A5���=�i�|����!b�b�s�X���V,�(ڢ��'���5�>h�42�q��
-��w�r�g(0E���n����K4Q4~g���l�� a�1�e�XHD�`#�=959��4s��7�a0�����D�0��:"��y;D��	��B���p����0v7B�8k��e�#܈���K4 �{�
 �m���5'��H/�V���A� ��׮Q!5��8h��J��u�Þ�E�;�'_�T��@;���ח��U��5foHj�D���	0G�}$��\��=b    IDATG�ߟ1mz��{���������T�p���^��S�*�����z�2��6~�Tki�h�}Yo�B�x�O����H�T��Q�z��#��"�e@ԗ(4YF(6��Z�`Ǐ�����ܹ�:vX:�r��YҦO�iny�-Z��b�����/~�KFU"�Fz���?ra7B�b�@��@s������:�?g�d{h�`'O��G:�6q�T�>m���0�
� �qڢՉ{�@�9d ����w~�@�8��� p�1�f��gpͬ}�>{�G�����U�9�N��Œ�u"g���x��*U"�ʶh��={�����5���c�U��o��Vki��I���p��Y �Z᪀. �Q�A��{r��	r� ��L��;L�� �ѦBݓfP"bEEf1���y��Qr��/͔�� >�q�L|r-7���C# ̱$�=������N4"< |�|��)��%�M��~��pX�V���yf��1��x��rҨ����s�8\W&�0峚	)-eq�Q�_�蜨�XV��Y~}G�CV\0�0	Y.<{��s�����P��7�v<Q���36ab�ūeKg���L�<O�P*ٔi���/���4��>�XҊ����T"��n�5��jj����'c�p�����|D��(�2��o�iӧXKK�u�:aǎ���9y��Ek���lμ��L|���;v�W��ekko�Ʀ��p����+F,�������F�m��������
[�t���9-^E����꤀S��O#Z�*5ʉ���&�Xt�.g`А(���녺�.p y��H��fO>��>��V�D�f2�Gi"���\���{к{�Pn�g�3g�͙=}��	��4���Bp�]]�|��PG�k�dx�MJ�����? bM �p��������NT��ׅ���a�p1.���4l~b����.f6�:V �6��pFx`�Y�ϸ� �p����j��u$�@���s*�-���`a<<'�\�
Q_�����-%�ː=��QA8��9a��o9��KQ�;�ы�����×����t~2�*�w&�"�)?�׿�w��`���'F�[J���p ���,
�u�{3f̪w�:s=��\�ٚU�m�U�<x��$Z��^7a�]��_�^M�c��A��),2�����@_���;�|=�?�>�x�;˺D��x֐u�|�+��+�!(����l��M[[�z�Fj��FX�߼�۱�I����G�p���)��;+�}Fn悃,t��@�ĭ��j�9k�4��.��6n\ocƵ���d/c��'�w�s�k�Q�5�Iy��k��B:|0�OM��W��8sB=���u}��V��;~f'�z;G��	�DXa2����~���!��@ uP��ϡ�H�l^�3P&���}�k_qpE�E��	��xf��d0��M����{�s���3��X U ��2P$� n~"��_���9��\��.L�Do0� >Z5c"��sPX ��'z�g����7�@p���\!w�5�8�@�E�>'���Rh����>� �b`��;�[�M�	��H/�.�0@��v�sF�xi�cBԌ�'��Ⱥ�x�τP�rGi��>e,������ʘk���sO���@��B���I{e(D�?�$�,
B�4iJ��^�?�N��n��ev�5���Z*�L"c�r��u]�w6v��Z��� F!�Y:�`U��jN�p^?����A��NJFdh��V2�{��nͣ,){P��]�K�㖑Q��]I?X1w~�N;x�@(��sX��b���j�Z�2i�gea���8R�#����K�ZM��%�Ny	 b�d?y�7���{,]o����,8��& ���������h��f`S����7Ra7�:�&>}�����FS���������?��T�
�!�J:��q�9G+��a'�u��� �E��3*MV5  ��\xm �a�E����y�&��� ���=�@�= D�����YE�p-�V��=s��m�{@�0���	���,kD�Q2�@�]����@P��C �yc�h�(? !��"���hrMb��h�0i�\��M"�9�惤D%�y< s�P&"�u�>\ۭ�tz����9o��~/�c����S�eNX�B�����J��ҳ�I � Z�5�%��q�?�f.���[�������X������R5�i+T����-8υ���i�BD�"�����7�)��66X���^����U��^�0?��^��b��;��Y�g��:8�<�´������Dw��U�EK%C2�sWü��[�ʒ����C<�)�t}ʋ��J)$	ł��� ��kj�;:,J:�	p���x�l���z�'k�U�������$�z̳�?��R��d����;R� ��4s�8
�s�eL�P���b�n�*iH�N �h��zդgNWϼ�.�Xڧ�4F��84�����gĽ2~Ơh �3�7��6�h�pW��r�	+��9S�-�仌��Sa��}$�枊����O8a,H����9�F)���h?��C�� �&;���yQq!���^e}��e���~��{�}�s/|-�e�K��B`" �h7o?�:%X��	+,�#�	�G`�Z`/Θ>�����!bi(��鞵5+��u�\9Jz�k"��է��isl���ij���B�l�J���S�롞��>p��Y���&R)+�r�V�/��5V������"��(b�>7D#y�!�h�4��M��j}\X�����b�����}����
fR�%;���j{��zCo���A
>��,H����^r�Ձ֏���D��P�#��'�[>4OBBh�7O�<�����{n��y��r�R�c���p��u�k���g�?��q��(ِ��IA���<��m��1f7��|q�q�r^lz�I�աW��(��p99��:5�L9�&����j��:�-�V��Ys>/�Ut
ϫ{i��$%����D"m�46�����N}nDo(�����XO��G�W���}�;4Hi�DXae<���^��1 HZXS�?�+�Nܓy��}�53��דlV ����ʇ`]��_���,�:8ЙX}�M��O�0Ux(�+����^�2�X�X�Z(�i�C�W�����ﭽ��~���v�4ѨkV)V��e�-Y��2c=��.^iώ�z
����	sa���ߛ��S��\�W�d͘/�rg:���9��N���+8X ^&\��H4�Z�{^<h>�P���(�;��=�L�� u͟�^�����Hl0�������F�_�%^��A��g8DD�l��B��Y" ������ 	������w���Y��S�*a��G��͜5���B�؀����w� /LH�=���V4:>�Ӕ�D�h�p�p4H9���B��h)�(� 0��VH"��eP&h�P9�Q�T��{P2h�h�P��JEà���g���c� Uċ(\?��c��l8kq�)����$��1C��S���U/��% �B@�F�Eĥ�S_��9�/�{(�ZV�@_�������#掝�����_[*�v|��I��E/r��ń��9��<?Bp0��r(i��ի9�%��4�	Ʌ�S�5�2��$�h0�/�!�G�k!�
-���Â?�/��Y.{�6mZn7� _��&�*��]a��-�l�l���Rҙ��U"D�Q�Y�����ł��
)4n�+�����S�J~]��{�H[]���[ �
_E�Rb����>�����3k��^v?��CæB�?U�L:���o�����$V]�ߞ���۝�� &�qSۣ��{��1���y
��Ъ�{�d�VJ�`:�����'�!�\
�Ā>�ihy2>��������"�	�c���w�#4X��8�8`|0g 	�K2���g�Q:T�D��!L��Ǣ"j&Q7X]|W���h� �N�(�%�b�B���1_�7@d�h��;�	�?�G\�U�q){��8]��'m�>J$����hd�?���_�h�]����O*�27�?J/�$��o��{q��g�x�R��pt{�{�A��G2�`f.��TL?���Ǉ�~�~.��%N^Ԣ�!/���b.�k(I���6uZ��sZ�W�o��C���/jum��/���J�d�r���/�CQ�������k�p����`�>)/�m��� {�hG�Z(��K�'�Gđ�9$1h�`�����?�_q����t��ax�B�Y��/
8/S�τ$�@w�0(��
�BY4`�)�C�Aw��������А��0�5F���@"̀��y܎�g�r�A�fko��K��J:W-4s��l4�_�9��V}�e��1���o�fO�����I�*��.��E2�J@��U�	`��4����@  ���P�8 �d Ѐ�*��|�*Aa5����c�!��.�
����3s-��  
�@�po��8H8�X/�<'U������/�3�����%? �$�ƺ#���!�g]�2UrӾ������lf�q
������Z.�����!�%��ĺ!�A+A%`�ܱ�]�/���|=��L����^w�y�3��ZN��
�cF0c�!DP0X;	��t����N���ok�.q�'Uݮ*��
��ҍ�_�zMj�s���רµ�C�p�cu��c%Z(�U��:�pܑ�߱�V��7f	�r��C�Qh(Q�N&�5pf�0Bԋ�&O��t�nݶ���==�?#�ӭǝ�1��s���>8xc!
Ӌ`�D�������%�@��()�;� ��h<����9|)���1^���v��n;y�Ò�rp�Vj�H5Y[�Q�羇O�%��?}����f�h�`0�n�r�cf^���ޅ  �s -<?`Kr?q ��7MH�͠�-��`B� ����E�>?4��5 }�w��� �.s!�8�l���z�j   �3r����h�|������R ��x&ƅ3ap	 �e H?����H��b P�)!�b2>r>��u����c8w����A���Љ��n!q}�A�s(�J��Y��,XM>������M����S�3{��W��khl�<ւ����{���G�����SXŬ#g��V��8�6p'�+��Wm�t"n�j�V�Z�߄�-��Y�Hᴄ5��n���Vs���Eע`����{0;��\{�gF���r�d[�l�$?��9�Bs�$�%�	qbSB���P\���$!�⊻-K��fT�h$M߳�>���=�myfd$�����5�=_���y�zֳ���փ���V�T�-TCX���gT�O��H �;FX���k��]r�O-�/"6 ���Q=����ܲ��==ݿ=2�G:��+�y�j���@�x$��[�lSo��2�'+�>�>��8m�U���ΟI0j�7V�C�vX{�~��=f��R*V),�Գ���n���������o�h1��gW��@ �D���-�' �{>t���j�i&�B��` �X�o�� ���%`�#��^2� �=��my6� ��� e (�}��z��K�P  ǳ�;W ���� ذL�2ѯciC}@��?1�U�eL� 	m�c�i�6�jG*.Yi���:�����^oL�PY�˟g�j�Pb��.�ω�	�b��b���al�� zyg,*�w������챋6m�׿�j_t�&j4�+��Ip�X�;�U�s��Ρ5��zO�w�����b�}y�x]��9��G4��iy��3��ʝ�Z֊�-\��.^�ROh�z�c�< ��w�>��	1�x�p`~�+��@��lO W�cx�����%@����޳����0'��6}�uw�z��O����G]S����+7o�FOo�F,d^��C���A��� �Z�c!1f�R�Z&I��t�^�SBQJ}���A"��5X ,e�q�'�`��g���^��XC�E*��G�7��]?��r��54R
~v��uf�
`F��k��ď>��SX� )�\�pŽ1��$��X�����R�@W���X�⻙����o �����Yx�G�`����c����B8�TAE<--tx,&PB����|���|��=��k��N:�X�B'�����bժt�(=��(2�O~	%��p�\�!��}��]�Prܧ,�����m�\ v����x2�#o��1�Yp��x�|�G��:V1��vIlǥ����546:��x���L��њc��1�v�{��Xg�#��! E�ܹ�O��}��O)f#��_�ފ�~�t:k�r��_J6n�$��%�Y�P���x���\�Q��$fG�/������|�j�:v�0j&�l�H��w��H-;�~Ľ��/`M�'#�y�hL����4�O	V����O`T�g��C�\(\�B!��{�sN�v�MwW,M�5��bV.Pf��_���f�^>/+¥m(��J�*H'~�c`�B[ <E/&wb�v�c((D��'�T��6s��`����G���~�|�q�>Fk"\I�y�Y���>:�x�G��������P��{Խ���s�9@u�X�܋��`�K������<;�����m$���`���^������ه�� &��]��K����]`aSo ��V����X�ܧ�`5����R}�����|�uJɽH�X|����"��y<�2�B��NUD��2:(+!�G&�;�
���/�Z���b��Y�y�P~|�u ̞��N�9�'xx%ހ��g�������ؑa͢������~g�w�9��g�s^΅7�K�ϙ�	�ּr�	ڧųy-V���,��kVZ"R�����K����[��l��(�� ��k�A2�����Ywoh�ٟ�YC*���?�Y����ƻ�~��+X�q��T�b����p9���?��;��1���>�Bry���UJ�S����ӯ���ۿq�Y���>f>��������I��Ix����CB
3�$��E��
�(Z�e�B���=�����h�W���p�'Mg�Jɚ���)cbx�-���v��[gW�����q�6f͜�Kny����Ț�Z�p]!X���y2���r?�G� �~��@�y"���z��"��ZM�	�D$�H�TJ4��$��p�s��¦������R�<�)�NV>����<₹GY{R�pn%�q/Ҷ�K��O%��̉�p���xMx)xP��TO���[��?��g��X��t�L�����c��b}:��#q�Jc�w}��>|/�������,�Jy5U�Z����� ����dB�(�J�8xW���+?���*��s�8~����=�W���6yJ��k�>��@\�x}���{m _�δP�d�¼L�k#�u����.������7_�ޗޫ�5׍���Ҽ����Պ��q��/���C"#�9*5�ϱ25�*~̐�w"?`���c��vr1eAk�c��p��sw=�t2�I�:���e"���y���
*k���$9�8MMf�����V���aY���:X̎v���V+��Y�Z�bs��O0y܄�6P(Z#�,zXT��/�ksg��C��h��`�t�LƯ�������
P��1 ���Ƶ�>���'H�*�zЕ�㗼)q٢K4Yd-�2Q� xn���6r���i��z�N�,�kl�V�����{l+jMV��1����_sl�A��������D�������Ρ�J\ �
�'����*��#N�	����,f���pn-bl/���#!�/�E�k�Vc;t�X��˟�2�C�"���7׌5;�F<K��<*�w$�oȦ-_豄ap�,����2����%2Y�4�;����N�����U+�iCRk��ݻ���@��\�x�I    IDATt�E��>��Ϻ�#��K��]=�%.�-�m��ܠQ�o���E_�~P���m�q0���ij�X$�6�yG�Dj�k�{�m�Y���}"0�e�9h��e˫��=�iC�,/�� ����yйm�|� ���-�1x .Y��r�ha�� ���@�i�X����n--��ˤ=��#.Q��g�Z����{i2�I�d���ϛm"Ji$��m���+� ��T)�p<Y��U!�wՕ��U�&�����_]� �_�qh����\T���������-eYr�L��D5Z��S�|��k�z�K+s/J���U���[�eK֠�x- <S��v�8�<C DupD;r-��� d@��>X������N��I8�Ȇ�������u�ߺ�)���ϖ�П���w�x�AV���<h3f�t�b-��L-Z\;�t�p��"������}�!�����G�8O�:#J��,��v�U=�.�i+V,0�-���܍��GgL�n���ם�)�B��x���/�r���h����-�_�ީ�o��g�3�����_≃��/hl8��lC:�S��J��?z����$>��9�*������?�Ο`�T�o �믻��]�B��\���bu�o�ץvP��;d�q�A�z��]�jչN��8TO�>��q��yˮY��Cf�iY�X������c�w?�%����)ƶ��_J.D�aGfB*8�X�ҭ;���{����e�>D��,]�O&e-^�ʗ�{�uC UqY�ҀkR`�����5�-��N �`. �w�EO�k$�C�9��L.��J�d�s<b$��4��c��*�>x����y(%���Ȋ��X����5h�g�q�d�s\���E��hav�2R��χ*��Q򉡼�
��=���r���=���s�<�V�ȸN&��HB��3����1u�+��s���i�?�i�S�Ѕ��r��p�5�x.	���)�0<��S�k���Vڅ�s��{�� �$V�Ž�������K�a�W�������@<�"���&��1�������[�t�0����cbC����pA����d���t���93��<���E�u�ڈqv׏dw��c���b2u�4��?��$y�V�b���NϘ6�9t&���|�2���O����x89
�o-Ł���y�L�@��Ǫ"�&:���@B��A���B�`;w�ԺzY�B����>�����ms���^�9�o�J��}O��W,d��:�Fp�[Z��D:��2�wJ2 �h�YXP��FÄF�$���Ft饗xP���}��>� n0�8X$ @*Or,�E�)E���J�.��a2�h��"�Ċ�o�&19�2��*��;�����-�<=p������Ce�M��Y9/|0E�xތ��	 �x�я�t5Ǉ.Q|����F &c�w�@8cL���`�h��x�=��� �\Ƕ���R�s�����B��9��do ˟�� 7Ή��kg_��k"������c�?��յ"ϲ~���=�l�?b�;рıh�T_ۇX��z�{m��e��5���v�o��J5n�R�Ə�l6n�r%�u~��{�0�w�g`���_��7���j�f�t�����"��2��x�4|g?1��1����@��qD:s���y��<[�>�e2$�%����=_��sx�!X>f��N���@�	N�>���o��V�<�]�|�߶m�x�>;���z��2$-�M�.����3s�"SU|6���4�L8L\H2 ���f�Q�< �Ԯ^�[��b�wv�ֶ�V��F�5_�5��%�wo�=��v��F��h���7o�!۱�h��y���C\�	�\'���@� 90�lQ��< ���H��&�{��# �dâ�\,,,"�+��)��YЋcb9�|Ѣ�3�X�XX)�`Cͱ� �(^H b�}�+Ã�<o
�2Ӹ~����ɽ��&.��<�7����ޟ㑸�+ә�)S ೨�����=� �����G��F���2�E3��L���ճc�O��O�y>��V ���?���?���YE�?��sƻ�9S��g�"I5 �3�(����wd� ���q����T<ԓ��k���˸`Fyĵ����YWح�����X�V����;$�H�$%�B�����l��ɶp�
Kgm0_v#�󧼇u���4��9d/O�1������w�B�\�2.	N���sc�+��{���x�믶���pgg{�=�����S[���7j����k���um��3�Z�y�����{DQ����=}u�[F��|�)�b�6n<�^�ZR�y�kn�k=|���U����)���Ҩ;oG���ŗ\��\}���I��Z�b�P���L�s�� �﬉	0a%���j�hR��ԋU,?pܞ����
��Ɇ�Ka��UϿb�X�-�P��U�f�(�P��)H��|Os��

���ʱԙ�ߋ�@����ŁkYu�yVX�,�,xz������aq� K��,(���� ��U�p�u�Pٖ�3�Ylx)�6,8�EZ��]�=ۯ
	���\�!����,"\ 1�����0tV4�b��d	�+d�+נ��|�'��C]���b
Xq� sWO�{9�a�0f9.ϗ�Xt� �� c��v|xWlG�>j�o�y�8�Œ�(�8k.Ԃ%p�ߙW�'ȳH�����1�����_��������v�R۰�����K��l��6}�|�0~���|C�8/��s�_԰�+���}��N����*6y��B�x~����R���7�)��*��n��6��?j��6n|���Z��>5{�寰Y3�z����vo'�{S<��8�7����nX�����k^s���a�%beoܞ�Ĭ����=�2J�R
���{��y��b®������L,'��QCrԣ�k_�]@-�D �Ky��'�?n�Z��F&`��e��n���\*����=d�����w0wsm���,(�H��������d�2��` hi���bun�`u�`�tx�,�,?��9�� �����>@V�,,HJG�i`U1��o��(րE�D0��(�@k��%p?瞻�3}ѕ�;�Z���k`q���Y�w}V�g�ǀ��҅��?���y�O�p�Tw�= ��
� �Kޢ���G��R*	L�N�g$�'�<��}d]C�K��s���ȣ�X�޹>���'�%ZJq����}�x(|`����y�#.�{Q@�,�������3�k#�>��_���y���J��n՘M�:�V�y�������c晐��F!�9i�|Ǽ��_}��LG��l�Θ�)p/�:�Zq<��^���&����֪��m�Σ���v�Z;�d���Eڑ�.+C2��|�M�8�b�?����n��.=WŉN��>�7s!����N9���=�o�tܲ��v��mͪ������u;ׇ
������:�TN���.���_�T8@�)`	������2�\l,?TG�v�$��W� �Wy��
�Ճ�J�j�׬��նm}�ʕ�gf���}�?��J����"/��?�#����\3Vu6��4�@������p\,y����m��� :�29��������"l <�?�����e�1�U�sJX� @̢�����n�kp��_q����{-N�3�[���11���\/ �W�g�f%� �b��xlâ(�7V?�f��9.�ͳe��&2��3U��.�lx7�[ �Y����<S��8d9��c9��J��$�,2�I-��s�/�c�O%τg�"ʹ�r@�f�xx�.��=��5��X$��)��:��Q���@
,�ݜ����;Pw���\�qKe�֬Yj/8�b������N�l���h�:+�Vȗ���?���{Tq4zG�I�P�ǎw�_�t��� �����^�;�`Jf��k�^�f�C��'�s��J���wYC֬�1c��^�� �:�I۵��i;x�î��[v��K,�����[n��C��zE`=tZ����C��>Κ1����m�R�;c����.�� Q�:��A����~;x��
Ť=^��3�z�D& /k_*^
r9^:�@%K +x��+\Ѡ@�`�:`r�^Փ��[��X��a{wo�d*XU�.����'�)���ޖrΜ�/��~��w�&^�g���w�4LN�^Ԅ�f�� � 7 �}�Sn�����-]�@��W2S�K9�&�hY�R�̤��z?��z�����-����{��e��j{ (1N��Иj��9�ԓ�e;%[j�^χ�=�
���?��8���zO����;������ ���H;B����kd_�)T(q � �Y�J��}���x��w�޾�6]|��Gx'�>X<�b�|����g5����jW4u;�x{Jv`1�	P&��P���%s��;)�����Jm�V�^b�?�;y�����'m���6k�Y�m�b�A�Ū'|�H���Z����j�x�c7�ڇ�>u�L����s��0�0Jx&�R��ϒD�K:l����lŊy6u�$�����BE�*I�q����=��6�i�����u����.>p�e��[ Nk�߼e�{z�Ӏ�1d=ׂ�ꬕ+�k�bM�������wϝ�i]�r�==]��SM�u��:b�r�����.r��������I�t�r*2��v�%�A��h��i"^�R��v�x̺��z	
� Z����t6z�Vk�h�"�3w�s��:��_)� ���I�A�,T~�"����lϳ�X!�: ��.e@*�\���\+�	@5����� �&%?9�~��nط~A�5�'p�3Wb��Zt�VO���X�ܯ��h��4.��K�(J�d�k�X
 �3���g�������pmx-����XR���Y�Q9�!��>ʑP�-4���1c��9'@�5J��R@����� 8cZ���?~�����&��H��Ϙ,
����h���N^��_��=p�,��VZ2�j_�z<&N�yα	�g: �C.	��D��D�% �?�2	�֗��dhlø#���Ž��c�|b���!����c�����b^��ҙ��ݷ��w�_*F�J���iu�����U��� %�@�홝;�ٌd�������_���~$�'��@]�t���~�*�A��;f���U���-�(��C�^��C��y���Z�Z���g����6zEJ&�� "V�^:?���I�$���䤙|���0A�(�������jǏ���������K��V�V2�4��t$�t�Yͻ�-��_��{*��k�v�zB�Aq���J��W� ��7�&)��ǩ�(IJܴ&���kW�W�e(p�'V1ϟg+�M��.���7ā�� �R�7�=��^ �u ���s~�'���iw}����u���&�/%�AaQ�=q��C��/���
���g�;��' U�`�B�Op�hX\�<���Pw,4,.3����q-HCG��Y���P2caN��;���KGa{��?���\7�� ��{�_�����i��Ӟ�5`��.�u�V���Z0�bi7q�e'Z63��.\l�Dƻy�H��:�hL��;��En��a����~���Q��������;O�4����-����]v׿��F&����{�b��Z�P���n���$;�v��{�?�J$�r@/�ݿo��3#����~�-'��t��9:�G2���'؟��y-�L&fw��5[��L����4�Vн�VM[_o�Z[�Y_�:��v���}5g��+c!��y�v���p�X����#L�%˖�%Ǥ����'���k��y�+���[��m��K�,c��7j�qaSm��N���G��)� �Zd���hI^Rp=^_<�:�Q�A�l .�τUr��tU?���J}kC�� 3�����A0y�K �v��n���@&zH�E.�ߎ��f{BD��[y&m�L���ST	���y�,�sX d��3����8�8}QW�^-,</>���#cDIO�PP�= ��P=�G�t�{#hK��uk�V�<<��<c/}��\����ze��3�ga�������o�UW��v ��?ng�\��@_�_������PG���3�S�$ׅ���_F�F����?j�dS1/�p����a��V)S�'��3$<��Kem\�D�p�ž ���&"����X�c4��'<N��/�ߺ��.@`� �g<d�~%��%:`�C�}�uw���i�N��q	g�}��/=a[��D�юu�lٲ���o|�Wm?��ϲ�H�s�� <�
�}N[��rOo�5#Y���2Y������k�s���-�(Y>�c�����e���LZ{�1k9�a���]�~�Ox&�*�r� �,� V��) ų���z�5��f"�J�+`�`%ԫ}F��#͖��,�1��u��ke�;����;N��e��/=|�J��fd�g��A�@8��]���� `���}q,I�ا�W��z�XT�J7��?E��L$a���(��}�p���H��[uQ�e-(|�8�hyql�~,`��⟵���!�h��`�����t�1��la�S��\��L��3Bm�3c�I1r�w<L�	),V+�`qs�LxD��.q�ߑ�@����}<+%)�W"�}��@��(����9�#��|���'�u�E��	�s�:?Q\1WD�`(��G�?���p��IXn��6n<�.8��}.�z&�]��U�)ˤ�s�Eό�{�^껇�����n�����qp�����]>G%&��ȳ��"�Q���=r��j%o�>m���HV����/b�4%-kv�h�5h��#���׽��]�֟ŝw��^�H�^������vǭw|����O��F������s�J{ӛ�h�j�*ł5��}{wz5O:��=�#��r�j=}�6}�"������PP�0�Eo����pR��A��2q�wדg��T\B$�N�T����	���
Sg春�p�Tm+�O&	�M�&[��#�u�;ޝ�Z?��f۲���*.$����җ�4��s/Ǿ��<���Tő��JR\���x,I,�ƢW�5��Q������U�< �X�Pyj�V��%/�-���5�/����i.spc,�47��.�l�_5� @Q5���m��F=D�`�J�����򈤢��&�a�g������έ��/����L��e��\���[s�7;�Y:��{��)��Z>_��	�-��X��={f�{�Y����<��cV�e0���e/}�{4ܣbP,N�w�������� 7�Z)X��xd�7EJ��
0x�i��K���k�T�]v�+���,���v�w=&�4~¨/�����?r'/+�X(���dMM��7�ٖ-[�u�a\�~j�g�>x��ʅA�t�B[�f�-;k�uu��D�7+�8I��ݨ�8���bB�
���:�k��+�í�:��y+7e���C��eqf�@Y@��i���5�B�xͥq����Ŋ:�c����_�Q Ɓ�J�~�,}��Jn+M��U}(Qr�)�p����+�l o��@ � B����j��n��nbN@�a�@7�v�;�AX�쫚F�2�M&�
}���L�;�ʊ����y*���o4�w�'��b1gMM	ה�� �{2���Ǜ9e�91h�Z�-j�`�s���Q��8S��jN�U����_��1<}�J��ŋ�Y�R���G�g�v��<J�'����Xn��]`��&o���Νv�Wi�EU��˿蜧5�o޲��{z^?���A���6A�3��3,��Oˁ����a�r��Qyoά�6k�\+US�8n�[Gdh�ؖ�@���ѷ�V  9'.9|,�����p��s�d+�7���ܼ���v��ak���L�EI�1c��+�c�e]�F!������ٳ�����\�,�_h���A���׌Sh@�PG0� l� �
Œ�Øb�3�P����L�|���Ǌ���)!��Ʊ��}�    IDATd��3( ��İ��U<�le<���ù�sa��	��"�˜!&�, �$u�D�wά���'(�V��8�}K&ʖL�l07�q�b��U�����d�r��ͯ�T��K(P��A8j��"������e����K�͛�h.�u���dA�3���빱p2�7����	�m��&��hs�Tow���y��p�*X �v�-c���_[{�W
�Li�<�Nk�r˕�����G��w�R��8m���nx�M�2q��T:�rp��8�b�W�����\+_�=q���FH~�}�IU>���KC�OQ����/�=��ּo��ckjL�@H)GFa�={ۮ����������,���&U����_�q�}d�364���+ �$hȮ`3c��R9 '���n�ɍ�N5�H������C����!@����>�+�CX��`�X�ϖ)ٹc���5�qCG�m)���I1?�@)fS�aQ]R�)����Ϝc�z����n��B�l���v��K�j�ު�bE =��gΘo���׽�s,Ny��d= �M�
�>G�����R�7_�V{٥���"o�k�:QAAeW�9�]_�}Ӧ��W��M�8ޚ��=������;�=��*�g���]{��-u���V��
ӧN{�i��9�埈k�I�Ʉ���7a�xzQ ŭ��D1Şsv׏�vK�~�,�X����[IxA�̠Ɗ���2�ؼp�1b��8J=�������ÛTSԍ��Ɔ�[X(V����~�����4�F�������w�������w4�7�lKD��ĪG#KRk�)����θ����PQ&v>jdþ,���>�O���� ���9�Z��k�W�q��^T�T�q��it�*����?�w�aI��
A�#`��QI�[�ϭ�Op7?�kk�[a�6��Ze�j�UJ9$<V��l��i�f���ן��x<.J>S��8�;��٧����3����߱��\ڍ����9F!:h6���ޕ��w������gKsY�	�%�Ugj�������:ފ2�k:ʍ��QhdS"�ͩ��
Or���x�R_�\�[xJ�����U���^�X�r5>�w��f����/�8~�%Q��!����~ ������]��Ԑ�d����Z�&O�a�w�;|���2^�%Ȃ��NYc���Ͽܽђ>@A� �C)�\X��we3��A��Po��Fߗ��#� f�U�o�Cy�Mݤ'�x������Ko�tz�H����]��M�<GEtǠ�%	I��E��C�t�2�z{{���O�
�# [Dȣ1�؎E�Le��� z5s)נG�����e�ןe]x��}������U�I+�)�7��n��-��>b��������K6��9-����ɖ-Y�^W�ҌA�*����爸$��y���z����&M��m���m���~�۾��t����à���{�0u���{�m_;y��:�o����a$ڇ��In�/���χ��^ld��ł�=n|hP�T��g���g�a�A��EF�/^8ٗL&0A3,;t�X|(%+�a8�?�붣GZWW��u
�T������.����>cV,T��3�r��NA�i��>�\�G���� ��3�c��&"��J�%H�$ aٓ�Ż���[(E�( zz����F���L#C���F���#m���,]�؟8���N����u���f��Xx�7d�/@!�9�^��zw�(ܛ��p���}�h�o���]�ܥ�I�?m˥�%��mʴ�6q�6u�l�x�Ű��U$�<W��p���_�B腲m�t�]w�[\�D�B�c��k����T]&)��d�޸=HxQ��B��,޾�^����8NC6����YG����X�V�O�>��;n���s>�=��ӨŇ�������+��O |�{h���Ui��cM�	�y�*�'����PJo{��<Y�	"����8zsg���K.۳w�l�ci��5ҵ+f�-�v���@�!��4v\R��5*�h�_,<�r��{V� �]C4���
P5R�0�@�` ���ᝳ?��{d�����V6��ˌ���Q�A�@]Я�r~���&su���A���m����!����9�z�=�}Y����#*U�^ݓ��|�袋�f.Á���s�]bm\�%�)�H�V:3�.>צ͜�u�JU�� �Hy"�'yEy,T�$�듟��Z���0���?�C�Kt��xv�R�@��˳�=`4��;������a1�ܳʐC�])�ĩa2\v�� ����Sq�/h�8��Fo�`�EE�"-���x�dM2y���O�#� ��=Ǻ��Ο	�d���YC*i�b�R�=vؚ�m��`�/T��7�������T,A�o-�nՓ�<��>�k��Ac�?i#�O�7��L����"D% �ÄfxY t�P<:�<	�m۷{�0�' ��l��>ۏ�}��ӄĵ��2����#���k�������V�^�F���G�g�>x&j��v2���`�?��J����͘�6��[��x�b���[��9w��SU/���x�Y�h�Z˗0�2f���d
'���)�h�nN�,��������k|��dqkjhp��8��uq�м,�F.�� 	��àO,h��GH<�>p�ӦO�����O���WC��?XQ-���>'�?�(E��cM��S�f@��M�H&��Vw&21QV0iFj�k)�,�IXS6fmͶw�V���9H`iii����r���' �MM������g�M�集
�R�@���ˇ�i�9��rI�b%3��� Q5O7�zD��*�xa�3V��?��%xw�I ��A�'��A��5r}���#g?U����b"��}@k@y��T
פ�o5�q��lq��^؍���f�zB���yk����˽��}@ۅ�δ�γB9$m�jP>)W�d���[�fNd}ui�O}�Ӯ�w=?%�*�ސ���l�G��u�<���,D;ɲ�1�^�e�{{z^7��_�h�jH��S��:�w���y�b��X`\`�9$e�äQ���n=�:&�Aޚ��{��J���"���J:?d���	�f.�梪 �<F���������󢪍� &F����82��� b��f���j�˂�*�e�Ŋ�q��1�����R�c��/-���5��kb��9�x
[�|�&F%�|��O�Խ����	>��I�+���E^F
s��(~W�!�9s��U�<�Ua�lM�[�֮4��:�SΘm˖o�L���-Rޝ���ۆ���%T,��{�ֶC�ٿ�,��bL<�P�d���r�(F#�&>G��O�8�� j!;�9Nw��;==��}a�����q��G-�ݯ�h�l3a�S���	,��ކ��U��D�z{�[_�u��Xww��#��-��v/�ݢf.���cD��⎁����5۠�/���2���]��ϻ5�A�hJy���Ϙ�8.��sw^���<	�r\��0�j����� {�(�r-c[Mdؗ�p�x'�cK�/V=�\��U�f?ߑ�����:ߋ#�~� �[��o�?��:Q��|�]x�9v���Z����x����>c�M�6߲��4N�B������s*����v��_}�
Q������K�+�K�bj�=*3S/�74���TOp��_��� �#�8,	ύ��~�Gp�Qd�);W�
c�KcA�Ť�����H=�X�i���f/�L[8�QjU�L������9m���#�왡�`T�v����?a�_=�cq׃?�E@I!ۡ��~�; %�q�ō���
Ń��lT�)���u�b1��(v���B�*�5J^T/�"�����!�W�R�;*�W)��Iu�D ��y~G�I��\�ߓ���������S6��a�
۰�\�T,���Ӻ�h�����V�m�}��P%���뱱Z�z�����?�s/��s�e$*�������Y��Kp��8��:y[���~M<�8#��u��~�7��O�	����?/��	�	��9y��M�ădo��*����:�8dmx�#}be��4:�V+)��l2d����0�Z��]���W�VP��?�\/]�����ON]�z�5M=�C숚0d�:hᡂX�
�dT�w��'?�I��_UQ�i�"�KZJ-@��2b|J�L�d�q��|Ϣ��,>��1�@U�gScP��XD���Ăǵ��S�d��x�������[����U+��mݚ��s��a"Q��W�	/�R��m℩v�K^扑P?(�<W���Я�q���J*��� ����<s� )|FYw=#�-C���Q^G0>��"8�;n����Qi��_��
�ؓ���xl����Rɪ�U ��B�8��� `��j��J�L��R��j%�V󖌺a�g2m�f�����l�R1���^�(8c���	�����>�B��,jh�C��G=�g\�DH��Ģ3�yM�9s�G?��� ��t��\��e؇r�xxT�e�����g�{�g(���8 ���F�-�	E�ꇅd0�?$v�����im����4�q��\gϜ�
�� �TUO���&V��m͹Km��gӧ�ɚ�g0���\��,Y��ZjF 8����[���|�;߶� �er����Ӟ�v�~G�GGY'�.�8��<�>����0����N�~�wo���O�濽���|�K�Ї(�@������Z[�ڑ�W���;��L��R�y�ZD���D3Ed�{�1 ?g�֘IX�4�HH�'R���ޢ=��6�Xƕ�R�-Yl�����Β�����&�#g�� /T6/�.�'W.�A�( ��Ή:��/2QJ%3�<}j�6���>�5��h��泟�ĳ�	�B���'@�<�*����8@�)>`�J��liJ?s�|��͟��,Z�9ǎ���-Y��ҍ��:	�C� ��c�P�͚��s��k ��j�����p�;k��P�V��,�t.��۝v�����~D��'��'���=P���l��[-z��x��>�/��)��܋�BA�u��[&��� �L����+7o�VOo���|�V��54f,ח�j�&��uM'3�
��i��fuB�����ِXLLJE��sTkE��+�<U*T��x�6����'��9f���V)�)`Ԝ�,W�)�,NF �A-n�.��s�vq�S|���:$9Tp���r�)J�׬d�_Mh�տ* F�H� �s��l���7Nd)��T^	�C�|�!���`��}��c�(���7��M�|�9�dYTH.���Ch�hu�W��NU攬��J��C�������?�����"+�������k�xUO,�Pճ��[�f?@���V)3��r������M�5T��S�[n��ٌ?��ɤ�ko�굽h����\�/u��� ���}�S���� ��5G<_.xŀr��� �΢LǼ��;�rȪU����`(I�ChH3�紶�GO�%��j^��R �d<e�]�R�;g͚��D�]R���b����� <���pl���冻����RkA&�5���C=�t"�T��;����l�\o�%1KE�Y��L���~���4�f�'l޼C5R�����I^����=�3������>��Ɉ�x�_}��սB%�i��JU�D*�ႊ/Z�e��y�O<���a�w��.6 Q�3���M�8��А�_)�d�B}�������F�-�xy�{�;$��PB� ��Y.�Г�8�k�
�˸Vj�qȠ`,O�:���s��	���P#��ڄ	Y;c�xKF�J�B��b%���[`/{��f�z�X
��q&�F����t� ���T&��	�x0ڔנX�EmK�Y�P�!es�Rq�l;�앎3fd�!���7`;w����l6m�R��r}��~#Nk�r˖Q���p��usή����y����'O����ϼ�C�����(����i���z�������D��FI^���5�k$��'|�l{vo��{�ZB�M9����T�|f�>{��m��M㖬��;g�-Z�0���b$����M�uY�xp��p�yNyB��ū�>/�	8������s��P�����ࣨDIe���ܵ���n鲅������;�UvA9c�����[�h$,S�%X�x��G>2T �kW�k;�:�Cc�{Q�,�(��w��]�HhA#>k�[�p~���퓌�N^_Tm��œ%[y�"[�z�{�rɒ� �4aǘ�4i�m��+㖈g��o2jd�blE��찏�|�{|�����k��z1�H
ʜ��G4\}�r	.��R���mΜ�^��Z-{��kjj
yh>X`����8�U(���T9*�=� ;����ͷ�t��i$�-jw'�Y*�����W��[:2�r��^%�h�;����O%A�ep�t�'�����A4iy�������+eȜ�J�����^�:.���������'��6�f� )��2��Fk9p���!���[&KY�͝7�� �.X5�s����������n�C�!X��5�d��A^4��;�6���+�:E����=`-�d���J��������c���a�(XI�h��D�W�,U;�Ia�����իz?�C�� �9�K,W΁�c:�V�7d�3�Pq>-Ķ��\%OX�Tϟ�>sf���z��r��֯[i]�֬�w�'�(�X� 64N��7\��o��P�Y�3��vx��ԧl0?���^L���8�X�'`�G4�(-l��+^��v�K/�d�R,dq����~2�T��=r=�rr���1=��\!gY�Y��?�W]��+��=o1�KE��)o�r��+�寸�z��z��c�;���O?��4M���sV���o�q&{���R��LQ;��XT
�s�Ԁ?�1Oaokuݶt�X������;P��С�ֲ�U���(nc�ۻ�m��O*M ��<���#p	�U���e�SٝJ�g0�z+d�X$FRA��x�3�:�S@ �PGG��h�W�,��� ��w��k��G=�K��:(�DUZ�	�sϪxn��f� :�?��O|���:������+�Я���b�@f���y�{���.��8 j%Ā?qU�9�S���D'�@�b��X�{�!����q[��L۸q�����W=�Z�ĬTIZ���I����.�rm?}|�ޛt�-�,�RZ�����+(m����K/���Z���ډͰp1Wd$�w��K.��z�o���J���ჶ{�km=d{����x�2[�t�-X�ĦN�IPK�����py���S���:�����v$�'��I��5kV�u׾��zl\cʛ��w��F�L��'��JO�\�
%���앶x�
�\H�ԜEY�L`$Ȑ���CC�[n�ś8��-o�^��eM`�SO��H�hW��9ܺϊ�ǭ����./�J5���mv���Ya��/���m��%6�l�Jb	��4�*p�:!����� rq喳���LX���G������f<�A�99�+��h
�!��{��?�f{G�, 	��$� x�y��\�V����Զ'}�R���BQ3$�\=��0d��/@H	
��P�;�g[>�}�˸b�q}����%m6c���|O�H�J%)��kk׮���W�%9+�l�3�-�Lv��3M6c�\,Z�`p,�^�i� ?���t�v�H{�;���hx)\���h��s�])�':�wB<d��q��gv��n��ͪEK7d�!��\>����	S�׮x�M�1�E���Wo��:;)�w*˿Z�>u���e���-�����s�H�IC��7�卶t�|ˤ��Ҽ�J圵j���nO��S"��.Y��{,W0L�;���>�$�Pޕ�����?��ݪbB�!�]�U|��x�r&&ނ,�z����h\�l"c�Z�b�۳o�:�-I]F�������m0t�( �9�C��e���^|-
�LLx\]^
�62��    IDAT)�~>��[^��ƌ�� 2H=�(� {���3^X��,7�|�?T,�_� cE�)�鱦q���0��Sr�cqn�	 �o.�.�?��<lG2�T;�6~�lG�K�$rn	*�RK��@�cɰ��Nr��^�YI^!˶��$��D���3g�V-�������Oٔ)Sfۜ�l��Y�;��К��\�`�����B���s}��G}�p�Ϛ��$Ç8���L(�{���X�R��Zﳖ�v����k�X�\�*�:��*��3`�J�~�^ms��̦bw|�{���ĩ��-�jq��iם�U=7o�bOo����}�M�b���7ؔIM�L���߿��\��K&:�<�-&D���6�׬�Xɮ���p�&����ʇ����qH�-��ʾ��/����E�B&�it�gܬ�kZ��l�� ]@��a���Y�<��Fk����1���@��X"fK�-�ӧX�B�PO|4�_*�MLZx]�E�� �	��k��?@C*�1�O �!���W�@�<C!z������\<���, �&���/�=���|q(��3��L�c����;��qh
�V�����".�^J5z�b���s}�A�ߡ��XCn�)����e��"2v$�4�<�-�)���騼�WC�
���r�f�2���s�F"d<��Y��L���<��-_��E�]���"�z�s�>������&���?q�,��' ��w�.��?�q��p�)X���m{�^K���>|�r�3 ���í�֟+��`ͮ��7m�y-��؃?}�n���!I�H#,j�~����+����{ð�O8�lz�2{���n�b�Y�h�����K.���B�k��:�&����m�uX�����}�h�
w�x�j��B3��Q3������2���Y|�!��1X̸��h� ���Qy�ᥞqK[��ʃ�M��%����`��R�X��w�p-��%K��i��Z�I$#�?��kf�cyj1�u� �[Dfn��H��ol��'��d|1f	��H.[� ��6xdu��c�d�m��$��.ՖȌe���� �l��N W	d=�U`��9����A�qY8(E���������op�d�K3Ͻ{eT�_����F��T�_�تs�؅���E�Vڂ%묯��|��QD�0�jV3J��	ć�|������
���44��ʜ��	p�k,d�Y ����v���k������w�[�l���h�-���<{��W�kw���nhN�6׮�������<������7�w�g%*p�G�X-��,^do���J9gG:�O���]t�:ˤc�ܼϺ����N5Z{{��,�h{���k/p���!���Sn!/��c1`v����,g^��s	(U��p�O%_��q)�{l_�6;ұכ��h41n���y���	�Ƭ\�[�Ry��5�KU�$����j-�&$�- �1��/n�I���ǳTޅ��#�@��ի�k �xW�?���G��]%�i!����'�!�?5�1t�E�w�=�`_��j��,V|ǘ��e�3 #���^ƍ(%�˼`�S������v;��ɤV)����K��ɂ�x3h�E��;�S*�J�l�������
R�[�\�_�xc �Z������#�g��'/�6�������@E<)��]��kw���v��sl�����������;h;w�l�dk=|�*��}�C��K|�o>c{�����ؕ�Y��)U.����J�~;��a��/�`/\g�B�;��	L��%����n���m��|�*��UW�}�{ߐBCV>3�f�r�X8X>߾�;���HT�� ���p2��|�FI�����юfk��g��#8U.��4Xs�ѡ�/��ր�,/ i�W��(	�[t~BC�09�������H#�?������L� `�2� fx}������E���w˾�U�vޥ�����{}�R�����'s��{?��@/�P �ԩ��`,b�
�]�{M!�
Y4���!�,����ˁNT�<��Py�(���o"^�b��֭;�6]��9�|+����ON�e�W�5�ĳKZ*�`�\�
v�P���'>����V�<ө7����@"��C���K�Ƶ1���b�o�������s�^lS�N����T��d!_��{Z�\IX�^�TR�я��������ܼ�KL(��>��l�o'��e�L�2�>��?�Rq�R���v�7l��U�y��փ^���?�tο����Ÿ�i9f�6]����kM@V�5�U7���7�n��@D�`yPPj��[Ա�57?cm���ԓ�.�(Y�"�Z$i;p��ԓ ����A�|*�'�%Ǌ��U@˟=E#���(����� �����qw>���ƫ�3�/e��r�ԱFh@���>���fl�p�, +`��z����?� �j�����[�@
G��)����˳y��}�f�6@kB�
�#��sqN5p�����4~J�gSc�����V�E�y�ԓ��J-m�M��i�d;���V(�,fiK$�<���ϸR�8������7W������%�Ur��ϝE<�tv���?�|�\k�fl���n8�����\�v��o�x֎w،Y���kǛ���:p��-��8O�����n��m�}���߾�ە�7���皑�>h�����h�_�-�?�j��=��}6�����`_xў�D���l9h�����]w]�����C�#���G��d��gR�s&�{��׹��-�?,(	8�H%���쩧���foW�M'���Ja��	z�v���<hǻ����=���z��8��8QG��:	�"Їw*�s#�`� :�Dy��~���=	EX�H/���*�ޱ�6�S d��R��&���]���O�'�:��O7.���E��wj5�1X$X��s P�]��(s���i�GM�J%cV��_{�'yŬ`U�7$wR�N��K_a�Z��unt�X��ڇ�\�Go��3qy.h x��_�5b)�7�����~N��G�w�0�bǺ�Q[T`qj=�i�]��~���k�`�7\�E�ܺ;��o<'�o�A�?}��n���[N?��r������e$��lX���]�Mv�k_k}�]� h�mmV*Z&s�����~/�0q����W�����V(E���o�;n6�~Ǫ�A�U�� �.#:a���z���E��re����b��sO!1e����b�<��-*b&̛� ��%�p�r�#���)��U����*E��$Y�����g�i8�
t�/�MI� �(�>@�"�o��+I^�Y$��*����0N����2FQ��v�w��E���)�E����N�`'�㆘eh<�c>@��!p^<%��1^��s�Z�	w,Q���Zb�֞c�t�*ł%��n��9e�6s�W�T+�ư�Qǅ�8���˾���9�so�L�ʰ�s�����S�#۰�bPʥ�#v��>��hsj���R%����H5X�T�;�Y2�`�����S�{ىo~�[�ӟ>4��)�v�������t�y$�@�/�\qk捿�z�3w�M�`--{m�Χ�ۭ��{(U�K�Y�m�s-�j�����N��Kd3 x�b�o�8��������@F�dU+<�QGh�^v�*�56em|R��%"���$���Y�N��Q�ki�|2|�zEQ�ꑤ��3��=�p����τ�?��Á?�*�1h��-����1E���0��'��z�� ٗE�W�I��%����3�n���߹�[N�`�(X,%��������@[��)��?�#��8��L���;�4*�2�K
�z;�9�ς���ȅ�&Mj��&{UO/�Xt*��05����T&�4Y���c�]In0���Ɛ����3���:���-���	�f���Rgh\6iG:Z�8���;�����^8C=�����%�^fM�B������/���	���- ���mw�z�WO?���>^ځ�?��^�y筱�_�?��?���zmǎ�]�s��O��d�̚� �R̃��H��%��ÝE����o}k��?�4z����?��?��L&ܠ�����?\�77�k��X�T�$��(Z��)�ʖ�d�>�%�F�^������j�Q����_��M�ZU%�>
62�Ƥ�?������v�n�±������^x?P����{
��E� +@�g�ƍC�d��J`c1�P�*���n���;h#�9 �𦼁<Z����������Ϙq��ba9C�2W 9�sB�: |����I%�CU�t*���>������:}W�%~=.�%K�yrd� �<�RԎ�gt��a��_�eμپ�>��%ܻ!��c�!ཽ���y�HZD=zĽ�'�|��Cpl�˯Y���=w�M�8œL)�����ǝ���t=aQ�$�1�$M
�8���T�/�d��f�&M�	��Z|����n��
�H�����>ॺ8r��ċb03�xXE�_�YX�d��
ϯ���`��m�3��b��~�R����
�Wl�S;�)�b��*D�����$��(�� I�	񏴃�B��`5�� {��6��O@�Z@Ř�l����h�js9o�5�v�\�9- �D�
�R��*�'ޞ�]��Ї>�/Zs>��Cm�c<��p�,
@ �x��P�?�$I�i�H�/c
��j$�
�k�܇J���Ϟ17�}�'qkkk?��1i��?g�$[�p�UJ�fR�P�͛�{����W���L�T�L���.X�Qt-�W�5&Bc�8��x2�B���/�`	�=�1O$��MQ���\�%j<�����$�
100�`WO�3�|X�K���7�s������-�e3Pqu	� {�ej��w:�,2q,fl+��Fݐ��=�)4�*U���X;z&��%����ޡV�];�c��<�Db
@R�/�g�a{��^���>��͎���9O����
p���ͽ��[�'���;T5��0��?���ͻ'Y D��0�G<3���w��|�� 8�� ˛y�1�'��Up�xrP�Gq<��}�W��@P���W�wE�n��ÜQ�"2��:��Mg@s�>G�mBL�RW�y8��k|�6h�Zf�_mF�R�X"��$ǁ���k�lm�Ԭ��B	�Z��嚢��2��_�����Qo�y}��/�o�>扏0���
/H
 ����3\��c`NJA�*�2Hهg�������JMwZ���-������Ƒ�J<�1Ȕ.���dnP&/������->�^kؓ��2�M�'��ŢW�� �%�TUO��F����3+ێg���P*��Y&��~�P���Q/�Lc5���._�$<Y��OF���k��^|X���\7�/W&E�d���y��7������ċ�nx��HOJ�y���&y%t%�_�+�|��R���U�Y'=� 0���1��X�(�THF��J�
Us�1$�Bu�6� |�L�W*��E�%�W}!�����چ,�����β��g�b>��wN���Ujq7�[{�7�
�@������y<^�Q,:<G����s���<&�8���Y��>�яz��W�A�<+B<8�����3��𼠿XP�����d�c�?
F�
�UISJ)%���jG��s*���ZH���AY�|��h�نA�W@�Z�u�	��*�'��Xaox���4�8ٵ;ةZWW���{z:��U:��������w�O�y��b��-^��fϙZ�UF���LV=i�%'T"�\�z�y��' �V�, ȭϺ�������"eч��pT�$8q (G@� c%�L>�ˈ#0�⃪�0��4�G���ƈ
�i�H&�W�.�"���o|�ϋ�EP`9]ŠU��/�|^�W�7��%�CUφlҊyJ�������Z]�>V1yz�O�4�Θ:�/^:y�)�q��>$-66f=��2����н��w�*j')9��j� �澸O����IU�ERυg� .�=F�:��^��H
���P��JӧN��4�z���K@%i#��˲R�h���|��>�C��,��n��i!�K�Ë��L�b�xSVw4�cB�`�H�y���\*�-V+Z__�<�ú�[-�E�@�Ѥ:�e?��a��H����-�g�fOwz(^K�j�s��X5xUp��&`�*�� դ?�e��A����eA,�n�
���$�D�;�� ���Bg����{�2/�`̊Ҕg��\΍�1������,M
����;D���3��x%|8��Ca�V�N^�U=U�٬X����t�rܪ��%bY�5�L�4y�54��L��
%4��~PBC�[Ro<ݛo�Kf�ӷ��Z�0i�'�a���H���ûG����_�Ǭ���L���^f��,m%~1�����j����������#�<|�i�Ղ ��� �@�`��~y���$��!@�Ń�G�n3����眀?n#�q��[�qo�ސa ����Xs�6��h������;CU�\�b� ��ϵ9s�[ie���*�~Z�4�����;��k��P>����C�/�%�幊g,�D����AF��V�!N����ƽ��Z�%ٔU�1D����ǖ�,�EsPF�"���b�x6m�<T�M�ζ
rj���=Q��,OEU=CI��4%ɻ��ϱ��?Ǫ����9�;g�^`����Tz�W�-�V$^���{�*������O9��
������|�	�X�h�U�n�h;C�.�AϙsS�D���/�N����2�O��W���)e��B�W�/\�.^�"��Lhd�������Y˒���-�4�xMx=h�D��;����IKO�[oO������>�S��w����'��b�x谵t�"�3w�U������g�
xVr�5����+��|�O�J>�
���>��{��� HW?��g��ƶ ���q���b�y����U�K��~
��#/�G�D�Z�W�2�D%�k�˜k����Hj29�P=�J)�}NJ:��a���a�ٖL�Ӄ�l�|�*�:s���d�s����H� ��<����3_[�a���}th�s}����
��QZ�1�Ƚ@�To�K�g�g�©F:||���UKގ�������M�z���?EwM���������{��]������ٚm)�R�Bh�iIDEE@D=��S�v��;˝�������"-	M@J	%=�������g~����g��eg7!	p�/^����Oy��y+
/?��4[nHic�nt]j'��Uf5��aM�N9�\@�� w:@l:!k������+�d ��;�c��L˺\�@��ƣ�-EG�Yˮ���?bd�U��D��W�o_��&��q�1P���������\9�����K��AZ�\RH��z�=�G�,;eq�:��\~<֛�#���La�tMi�^���w5�rƿ�y��|7��9�����!˘�ƌ0m�1���H��4Ǝ��c&��D7�`"���L���η.>�hU��c���+ĭ@�����r�����%4�����+��!���z�o�Ĺ���_�O�s���b��kim�����g��_B����
�� �ߵ�\ʙ�d�b^K�T�F͞��c0}���$0��Lw�:y�N��G � `qa�{'�/�+��ͨ�9�#�X�~��e�ǳV"�g=��7n����n��O�lZ/|~�����C7�+��G?F�<�2�Hu�J�R��7o�|��	�.��8q���-��;����m�ē��r���g2�T�Z:t��7�+�c왑6b7�Dp��(�,����� �����u�x���0�F` ��4-2���T�沎���5��w�)�OO���D���`�UW]�g��>����زy�ݻ�ݽ����Ne՘�葿Z'�@0
zy�Aq�V�Z�Jf,��9��Q8ɿ*��/�3�F�Ў����-��M�g�-r�PUgvЏ�3��S1�e:1c���1�D!��.�E�4"V݈��&6�    IDAT1�(+���l�p<��+s�y��i޹RKU����,k��x����R.������P�/5p|�n�zj����+-_�kZ���埓�HDҚ��f��ڠ�!��Kn�~�ݐÆ���m�J�}�D
ȧ�uTU7`��Mx��g���ΰ-]�ʍ�EC)9����R|>��[�v�]mh^��څ�
_��&Rq�T'`nݺ�������E6݁3'�S���O��"/�;}A�
Q�3E44�⤙���u�+M)�ƸX���mZ&�=͖^�[ɋ  *|����O�'�F�P<D��4�!�/�2�����|�L�S����ez	��wU�������_T�qoLA�C��XA��Cy�K�����|%kS�2	���g�ƭV�L��9�I�X�v�Pd�����ӳ�z����,�s�F�P�@߱#?�k�a��V����g��������i��=���'��O�fl�(0��3��"��aX�p+�"
�(3�`+��n$q1K��\�$�:ȏ�y�6V��4o5�SXB` �oni�~p��/���3jk-2oZ�I�B���r��l�
�޹�<_ח�Gn%	 Å�@/K�)������?�ً�h !���2�Y�C����6nي'�z��$Ba���p���1f�XdҎ(�ii,ء�G�
��:}h��v�Џi15*�����ػ7n�?ӧ��I��ǍǉӧXrD8��c*r��,�ٜz��5��+����c�f(ȇ�A��`v����H�6��x ^/^�{����'YR:KTV�>PПn�A����+e�w�V~6.,C�)3%�W1
�L4��*�#)�;p,3RE;��s"{��2�'p�e�_�p�u1�U��#�w��|���j$��رk7�T�Y�R`�Xv�:
�T�hXiL9��<��޹ۇt]lh�c�W?"!Ge�HvPkl���k�oτ@����$��#hjn@.������ѳ�s驝�Rɜ�|(���'];Ѩ#g����`��b?^��!JQ���tv5D�Λ�"W���4�
#p�e����"/i�^
N��i���J[J`e��xj�fJ��o���6y�
�tM�k�tHiJ�R���S)~��?)����N&��N�F�
WYos[�� �H!V"���#hjj���G�豣1��s0bD�-b�&�@G�������7~S`�����%1O�����r�e�oP>eA^��ٜ�1�Ҏn�����|��cu�ً�Q�8sYa[�q�- ���:
� � >�w�gT����}O�K�\b	�D��*{/�����`���x�����N��[
W&�᭭8��3��:�t��+-�i`X6L��u$n�D�P��ތ!	����{L�����a@�]]��gFO�˸ TU$�t�?\L)�"4o�SE:����k�{fΘn)r
R�`��,Z���v�!��"+��O��%�,K�x�����%ȿX阞�;R;��[�>�j��x�K�;�t�"38x��딿�wޏ�+��5��3��Vz�W_w��������RN��}l��4����Ǿ�ml�Ej�|�|i*Ϣާ�x�/���ۘ��|�����t��c<s{�g]�[��7��,�h�z�����wߋb!`����(��DCat'2�j����t�"�[�]��j�c����k��I�����5�� 8��;X<��q���G	���~N����>��!�����b�ݟE^�-�7J��܋L�t�����(䄾�k0m�q�1P�3��}o�ހM^���b-�T������|ģ��r�x}��e�9���(��ln���<�1�&q%���D����5�*�����{����ꫯ�s�������h-��4���f@2�s�������o,J>�6��������]>�t��b3�ѕ��3N�[=�'uD >��7(��u1h�̸#D�~��]3o~`�!��?l�� P(&m3�Ǎ&R1����#9ʡ�;��H#�A��n���Q�,��:�*<O�ŏb!_ dϗ�q���E����X�
pj����ek��Ϗ"��C�_4�y�	���2W�sW���S���Q��A�g��@��5*�2�.�r��vr�}�qN�
�f��h7?n�
șu����}d��d���B
���(�Jb�I
�5k��?]��_˥oz��t_ݟ�{��ʲeϛO���G��$`�u���<�����������u�7p�N�gL���^ U��woL�g��{Nq���8��_@??c�n��P���TWע;���K�3�i�%@K��>AG���5҃��?��������\����p���"��D0����²�F�le�y���	3����)S1|�([l�,�]�|�M
?�{��Pr����j��U%�O~�S��\ ��4P���'ٙ
*�i[���Ի`D~CUHrQ�r���]XR��~_+�+R+�
sA�cˋ�H&�6�Q�E�y f.8���,V/P0.j�N���Q��[��aaN��l��,'��;>��ʆ7��;>�}j����̆�.Y�
l6��X�h�)�%���6z(2�iS�dQ���&P��p�B��}���s��2�>���RiLl1�$`��������i��tPd!R>ւ�|V��/WcB���B1�N�0���=8ͱ�w���~nŜ�)�.�bP���kɕ�ci�X<���_����w�{�:��c	jn�l�*d�7��dZ5}Y�
���W�p̵_��A�We�]����u�x`*~׻�X���	��.{o(&�z ��^���fR���O௩�K9���w���a��عk��SScƏ���3N�~�������sK���O������:�ނy?��;n���,���8G�>��C���LC۲e�|�Q�;���0�����ο�ǉ3Nø�l�R@��G?*7s (35졇�x��i_�U>w�\9�L�,�O�� %�kA{ϯ�a5�8��6H�Ks����ٳվ��B*܆�a����5��!g-n �Ԇ��#	
�S{$�dm�>ט��:�l|SH r��M;��A;߹-r(�]@�.��.�Ի��&
�a�%����	rL�%�����/?r)���!�r-q|d�p,,�C?p0�xe
E
K�E�\|��ˢ�,�Hԏ|��K�_��~��s`��Y9� >Q�	U~���06W�sI:�Ɓ�E&�:�����
~�r�oB�ד
�s~ow������(���|�w�C�	�r-վ�/A!�GkQ�@�W�C��*��Ԟ�P9u�)Fa�����Q�����2�g�����g���n��I�Mwa붍xq�2�]�Y�c-��s�4kƑG���M�X]$���7��'�3}5��_0�����gZ��ITǪp���ٳ�J'��Վ�;6a�ڕ�XҜ%v����ޑDC����ך�g����g�d�YH3�.!���z �+'����ȇ��\���'��``��kj�Vֿ�x���M��9��,�ȣ������hf&����ȕ���g�,ɥ$�1A��1wF �l΁-�P0Rr�el3�	v��c	�sHf҈	�A��	������cڤ ��|�H0T�hx�Q d�����~ݿ$t|�����YՏ*ӈ�'��I�܉hU�	��6|���m�Fb�:��Y��C�e`�-����y}Z]�R�!��v���>��6�����|_�o�~:>G՜-�.����.}���o�G�����/o~(ʆ�xȚ���ۓ��������X�E�l
��*g�����4˂+Q�H����)�bj-���B��/�Ӂ��ͣ���ǐ�¢���g>��F�F��R5Y)Oz�����>S>?���5e>�B.G���ذn��چ*r�\&�5��b���v�L�s�F�Θ�/�+��)=Ͼ���1�����ߏw�o���S�rݼj����$��a4�U�ww�S��d"���6��&����۶�D2�Î])\r�[q�Ygوs�٨�����G$p���[���Z;"�Y ��w���hCie�@�/ ��UN����t����H�ՍƦZD��X~n�u����[�)u�+~�3��O],�@Е�s��s�s��;���Q����(Z��I'�� �pO�����\�֚�F��Ӊd"��a���]�W@�#Lh�K&��8] 4�0���sYz�z���6�;�C�lٺ�R[Z�͔D?���_&ldb<���	�g*�A$\���v�wU�0������%�3�``n!]
9���v���)�ڣ��khmѰ�P������u���;�mn5���F��b$�j�N���o��xI(Ïp��d�w�Ecc���e�0Ǎ�fKZ?���\�,�0v��_ l���xD�Ae%E)�Rp�n�Z?X�_�Ϸ��(��8��5Z4	>7��I'��/����g?kV�R��\<��<r�n��ғ�2��y�F��1���-�͛v"ѝFWg�]~f�<�((�)��寑+d�)B�m�q�n�_�����U_!h��Q�F�s�������v�0��S���ֶ��7�`��lټ�`5V�ۍ�Ǟ��~��f����]�(���G>�[lq�zR(�˿��� >����~��D*gn\o��P�}�9�����|s�<'�e�П�!�u>��[�@�B۷�㩿����{pͻ�j�'���R�r�_je��H����K�੿>�a��8��3Q[C��TbOp)�-L�n����~[6n�I�gb��1�{b_�B���{�X��R˪�d�YhF��T9�aAD����]���>�V��g�Css#�:�4C�
`�8�A:�3Mه4�LWdp�
�x��'�Pi⤣q���/cq(���A��OR� �q[ :;�x�'�Λ;��KY#ΏO!@߹��KMxؐ���������SO��L���5wV�*��P���}x~�Kv��SN��)cM ��a�@�IQ�_)S.��aǮ��랽����X<����8��	���o���;z?,����5F�C���s}�k_���>����Y�ϦM<�^����FMT��ɿ�c�D;���?b��ᨭ�F�Ƶ���0���JᕗW!k@[�5v>�w��^�;v첖�[�mvsPR�z5��_0�{������E��TL8f<>����V�Z�g��N<a��v�؆T�u��ՙD[�&���qL�|<>������I���B!S&ӹ����'�P0����C�Z���Be���J�/]��WҾ��M�.-���@��-"�9�~��Im�\6��/��IG �ڃb.m�j_>l�`A�b�B�y�`;vv��G�!���/��p��@�im�&�F�`�|h2S���kVo�#�=�au�p�[/E>w�}�8�R>f�d���?��#X���q��:�(�3=�{�=��.��L*��}��q\�΋P]4�`UU�4g��JUz�e_۷����?��#G��K�"_ �e-�)�r�&�g9dr��b@�����59n��v�t$��P`��#닙h08ZL�62�B��r���9gOGsK����Dssn�S*��*I>G�y�V�}ϟp�)'cƌL1��ǥ�z}�.5�M!�!��%�-�O<�3�:S���v H� A?_�b*�|ϴ��c��v,Z�8�	��yfS#�Z\����^% � �� +����-1� �����d	�%��#F��v�l��n^��L����-Ƨ����OE��?kּ�'�N�6MMðr�ˮ��AgWk�lB&�N|�����_Cu���.������+ʬ�ڻ�̟!���>Ǖ}��q���o4M�ޭ��Ow��9�M�ݲ��DW��#�Ύ֭k3�߰1�	��7-^��� ��M�� ����ċ;� � ��A�3!�23�߁}��\���Ո�ʄ���_�/�8��Y�8�� ��c<D���M�C0�3�~[�ua�%Ȥ�����Q��ȹwf:�e��4Sr�(׬m�c�=���:̟w1�$KrJ�����ӓF��j<��X�b5��9�?�l�U{�h�tG������,��YtttᲷ���z�I�O*�	�ְ���lX�>�c��/:��=�D�˅�D2�@$
�$�r�0��V<��X�v=��0	g�5��N��R�9b��~?��\���6�����~�aÚpڜ��:�� �RK��y�Ɲ��_1>�c6mڂ����8�sp��Lw�Ͼ/��K��{'��!�z,_�
�?��<�TL;a<ry���A��qə��4��wo
-z��.k=
��rZA�V��>�����Q�>�W�J%�����X)ۇ��~T�W�5�D��/Z[M�a;����wYV��X/�y�[�����N�3@W��5+���s��!d3�\��l ]�Y��E|埾�`�ʺ����?�굫LY�{�/�������@d���#F��|��e\��n��4�8 ����TPƢ����[�+D�qs��x
n��F����n/�2������6,\��x����9g��{�5��m�L+@���[�l���c�+8?�@)n�]���Z�3�8�=g6��X,�7��#�4ͬ�1�7RÆ�Y�ޓ£���T2��_~b�r�����ϥ�Q2߶T+^Y���|��:\�ˬ�]u. O͛�T
�]J��F��ú�m�5�$?}�{}�s'���'�s�JK>C|o����i\z�h���=�����/C6�|�e�h۰�-�*��r��"�NWe�u�.����g�o7���X��q�_�f.�c��|�k�1�KQ�b1��N��f:+5�?���w���0�1�r�-K�.'
�_v�"	 �>֮Y�|��~�N�Z��;����Rx�o�G�2�=�|�
K��h�������cǘ_��DP�G�>�y�|��?Sx���ٓ��E�ބ�e0��;�̨W����װ�����J�+�{*��
��J�KqM�'�?�f�2w�ҥK�eFk��t٩����i����	ذa�~�^�7�����/ K~.�zC�wc��G�c[5����'>���aX�n#~{�-�M���R��b�����A��e �`J�>������z��]x���8rT���]�{M������љ�捛�i��j/����5r�Pkb^��f�?>^y�#l���W��c�a��ٸ��������M �8L�
�-i�}��p���bx��U��3�.�ɓ�@0�u�UV.����o �?ņ�x�ѥ�z�;.B4l��������X�ڳӹ(~0E�P����.A(\�K.��/�p���L��.64<�ebVK��۫�x�_�~�F��'Ok���"M"/�P[_�\&��D���5�"�L��������s�%� VC-�Yg�nT�� ��a�0RE��*{��X���3;����ٵ˄K0A6�<�����ۑ�&QS]o.��x�<�֬^�Y��a��V���teutbյ��l7������*��;���=6�����OPW?��2�v�4����~��]���?`ƌ�s�$:��]�1���z�5$)+��T�a�O��4������ǌBw��(��6!���+�D��h�hG
�0v�N��+���E.�L(�]q_��G�sޥ��@�k�B��ʖ7[HnQ���������R;ŧ�=̿�׮]kץ��Һ�3�O}]�~�>�.��`ێ-�%M7�ջ�CX��{�ص���}�1���Z�v�e����^�=o��/5J3�|>\r�[p�y� �����e�b������2��>�5u���@ۖ����_�N���~��X掸��կb���fR�8����$��1����shp�H�e��.�/ҫ����`��-XH��gҤ1Ȧ]Jlk��6����G�Y��w�!W̠:V��;�X��Id3�u�y�U�H�hEZ��Z1z�K�?�^�;�	�PUU��k���Ï���W]�6�	�|Y�=b�}�Q�ݳq�F�m���mZT8T���[�5k�aΙ�b��#-x�L ��Mhmn�豣-��qs6nX_���~�b��O��@����CJ8A���    IDAT�������l��=;�m�f�X��b�Mx��'��P�K.���_,�b�w��13z��֯{�V�������I�m؄�'LŌ����k���c�����Ƙb�q����B(�@���������a�Y3��\gV�)�5c��񨮪Ǯ]۱e�Z���.�T�~�I1k��Y�`ֵ�y�9��˦����-��=Q��]V���Ą�c�򣻫Ú��6��@g�[�m�Ν��L'	נ=��,B<�,k�ƛS*D�AyU�W���ڂ��H����}����?|_i��!�s�e���[�j�^V��|��!�
N?�t�T�g:�n�Kصs��@���Hg3�ҫ�fV�K/�6���W����܉��.,\�PO�Y���P�oni��������1�A��uj����x�ϓ���ш�n� ���ȫ=��>�4^X��Ip"���>� N�}:&N>U�l����I+A�L�d03D���>6u��0b�H�[�� h@����ޟ\DFJ��~>ܜX�:m�����X��l���w�-s���I��M��L<u�����8ַ����]����)�w�"��_�֋�P��a��5b�䩨�kp�7�70f�<�ϊWV�i�}�jq��������Ǝ3�j��Tr�Y�ʺ��I�i�},��U�0��,;)[�"�ǔ��[u'��\N�֬Ya��-�:;�x聧lc�����\�8��駝�|�o�[ca�%��3O����m�_�����!�O�=Z�����Fw"oEl�\�����+m�؋a��Eذn=fΚ��'M7৛�����8�����b):�v#��Buu=~��[��쬳g�e�0d30�9u��o��@8��ӆ�<i�Z���W�5n���'L7Z�L>�qG���e�3Q�*ڸa-6o]i� �b/,{�=�8�;�\L�t����Ģ�8y*��u.���GWW�7;:��ol.|�l����c�1ۗ�1�_�ֳ��c�o��,)b^k��\KS�Y����T\��ϸ�<�v*�&����F��شq=�a	6mjC!�A�u�˙�Hkw���8��3�٦r�=��w��]�v�ǧ��?����"���l�5uHuw�8���p�EZ��ݝX��9�̙����S�Zpgډ3�3���n�����ؼys��YY���������"�b�Y��O�w���\D��SS؟�}��I*Me����ތ �s�������QG�1�3���N9���
w�옝ǚ�+L㣏���E�6��[�z	jc�( �#F�ńc�������*dy�]���=F����ex������dc˴A�-��`�6ړD%ScGb/���æI�U7�~���u�}�Id#�5���N2_��9f�6+W���V��Dx���gA̿�\��ģ"N:�TD���,hcЕDy��6�>��ۆ����g�Gĳi��@um���#�M�,_�ľ�Фe�K/c�ɳp�qS-B��ة���[���֬{ъ�BA����n�bU8�hh"wL#F�������+���M'���{v�et�btIΜ9�O8��+hI� qԨ#��A�H8�]�����9 ��^Y�Gys,�j2��4Z��q��i���?B.��/����L(�^��>�{v�j���z�`���_��_���Z�5n��3���֯ ��?�9ۧ�����I�?+������bP����n�E*k֬r�D��{��ZP��9s�c���1�-��H$q��oǣ�>�)�Km��A��@�@>��?v�����;�\ǟR*n!�15 ��ј-�Ԁ;w�4ʆ�^z��wS..��'L�����7e���5�QV
NБ/Q!�����ӹZ��)!3��4o��g��|s瞅Y3N,q��L�oji��ˏ��V%�k�V�?����Y�=�l=�HG��Bc�(TU�ώ���S(����c1m7�{���G�Ōf��u����BC�00W���8R(sh߻�,��K^�Ë�9���̓���n��I4Է���,1��Mw�5�hߍ��^k�I@۾5�+��#��3�c?u���kh1����WU��u[����2�}̽�|�9�]{m\he�@2�t�w�EZ��oCw�?��ο�0a�DTW� ��Y�OK�&�
E�2L�d�;en#V���;�c[.�w	F��6�U8X���ᨎ58�K��H,׍ή=�h��K/��SO=m�o޼y���2¶P���Z˰���u�T�,���N��)�w�h۸��c�%f�dShj�Z�2;���YDcUH&��s��3	�}���a�fd�yK�e�?W����wߌ#������Be�y}��3%RhP�E�u��FL�"�Db��(����V�y睇�有h�4�R�o7� �G���R>I���Ltw㩿>a�E,2WR�׸�J������7���OM"��t�3�	J�?�S�֙��,���0�E��1N	ݨ��}��f�o,�Rր5����rQ0����9MEf�9��/e��g���(��L�C�|&n
ˮ�pՕW����@w�����K>Q�.�?�����"���M��M7b��H���e�����;j�Q�2�̾����sK�����_8��0�����d-��M3E.gi�N�8Ͷ�{���m�މ�-Ɨ��O�h�oFu55_f� ��U�1��&�Gx��'��_�����U��,!�\��L��0��-%0_�r���
��w?��O8��Ӎ��2_��1�ч`�u�rM;�&���g?�)V�Y���w-&M9�h�K�D��'��j*(X��	��꘽c&�ړ#F� �l�s�C,,еBM<C-�� 
�<>���z�U��{fO�n�,��9��S���4r��ձ�(���o`��Mx���c��wOյ5�˰��DB��,��*�4���;��o�4Z#�DM(H�z��yy����ތ�5��M��%���ܫ���-���ζ�<���x.����*c��!Z�sΞ��g�RBp�%����?T���1�F��G{�^hB��6���"��ń[r�z�5���T�~��@.�\�}�J��Hu'��@��#�iy��H�B]��n�fA�%K��ɕo^t�ܨ��\X��9������^z)���
�F�lق���[#��G���V�'`k�_����T�.����@�wް����ry\~����>�qJ��aʣ�8�'�p���6[�KKK�}�{1bdS)>�F����N�s��r���x啗��}����y�7o�c�$�u5+����L�|2���p����w[�ͧ?��3
���8��
8*
Z�Jv�>�X˖?�[n��=i|�_G��<�d(�ppEZ�7[�TM����p�w��{�ԩ���>`<F2jst�T�/�\�b������ ���obÆux���o-6	�|_'����	���eEV�`���}�߬0�C� �Zb�V��#���F,G�P$%C�����L%3֓��ʀ廮yg	 E]"��3��T�Θ�
�mNw�܍y�.��g�m��9����UE1˭�.|�_0��B|?Ο���[kwO/�����@� �G�2)OR����`���c	�7\w=�=�XK���c���5��Y�O���B���U[[o�>y�dL�t&M�d������L�,e���|�)l޲�h������
sO��7���6s鳙��L�&��<S�"�*�U'�{���䗮.�<�6,w��=V���=��w��]��f�� �3������q�@�[�8�>��{�\^��3��mWX���9�b�JI�GkJ��|7f8�}p�u�YIw�l��Vk�n�Oƍ�ϲ����o��/�%��s�W}�@��>��������+�.�m��vwZ��EpV���Kˍ�+�̚�B���j�g̜%��	aG����\�Ɍ�p��Ԟ%�պ��b�����������1���q��e���]�������|�Q�Z]���C�z(�'Y���*3o�k��S�rt����OBC6N��Hi�^0�k�87]ݝ��׿n�T�gS�S��"�ý��<^~ �oޗA]���7�lV(Ӻ�}*��r�������q�l>}.�G����ɬu� ��i.g�K�?:W�cj���|�u�p����-U�
�mQ�g��"���MWcN�?��?`Ŋ��;0q�D|�S��2m�iS�I��r�G=L�mj.Ϋ�~��x���ֳ�y�6І��o|Ê\�r:z���p��ӜB�*�a��͂\��R߄J������c�Y����3�\ݻ�F��X����.!��\Ι�Ȕ�}�=����fw��ח����	Ǣ���^承���5�	��ZR%�/p�W��SL���8{�7���\s>yi��p��'�ۇ
�2U*���;�k��`3�>[~WIx����S���]��z���>��h^��Ũ�A��aP�B���O��O��3œn^
5�mR0+�G�}�kMy�0SkC�$כ�޵��$ �����n�����������p�X������<����޻��x9�,��O�Q:���X��O~?��O��SO�F�R���9ܸ�ٕ������fk���ݍ�����J�����GW"� �]�����C�5�����0p!�s�y��>�7�s��Z��2��k�E���6��s��eQ�gq75�)U��[g��q����,S榛n*[w^��2}J\�|>+7�O�Ss��M�Vp���y���l�|^*�&�k��XI��k��(tLP��Ҝ�7�T|f��_ti��#KV��+i��%�3��?�߁������@��>��WZ��?Z����g̭C�g̎���ts�QY���s��ˊ�Kq�
Y�"y�>�?�'&X��N�﷍�~�Cop�?4��c5��4�}ьg�We�X�/�R�����4N��J��1�!^��z\�W_��JD�'�A�K.
�?�;Ǉ���$p]{��S`���ečB<���E4�p"ë4 �ݧ)N���}�ƍ+��qC����H��y�	��ɭ�}n�� �����bޗ�?��,i���:+Ҳ��$���
��j�^W�B�"AR)�J๪ %�����r���T��S�j���eM�	{^�;��	׃,!��[�x��i��)P�Q��?;����˕ƹR�W
��k����ה�s|��x�	k�Ƚa�%>�]�F���ԓf�U~dux��!���h�aY =-��&m�m����F$['9��`�� B��w�X�e!�}��ɟo��?�ϟ`Lp��T�s��I2���N���DN�����G���l�C!z��� ;P7[������U_U�����X�?�~��_ۦ%��%����njC͟�d�,�� .2�ļ����PY�CAI��c���3��4Tj�^�qf��`�K�}��Oa���,��֟���1.fi=��~��aM�XZ���������{���l�e��ɱ&s's�Y��:��)��b�.!�w~�N�JH��Y��_�u�[��������i��X�g8���?�b�0��H>����%U/�MB��� �<=���^ӫ����ͮ�+�Y�\���,t��(��뀚i���$�q�8�Y%*��1��]�a,���{��/~Ѵ4�T��Wr2�-G��[���	qik�*cD�A�=5�z�i�H
��n.��el��.����O�����e9h2t7�閠��?��Σ�e@� F0�Ї>�Oo�Jc��p'��y�FL%Gn����z!�݀�g�u�i<^�Z=�i�󹔦���5ſq�8�|g�>�@�8	2�Ko7��u貚z ^kDs�U<��z���޷T�{��������������$ؗ�X���:�O_2����4.
Uj�	�<N��?hr�?�k�߻�}B��]���]�8��N	�D�f�]�L��ޚ?��c�l+1��tKP�_J�/95p�ɾ�8���ÏW���ڠ��㩽3�[�L#R����I��k��V��S�3�ր����o��4L��ILŀ<0������7O<����]և��g���g�	c+�w�
����TO�+��FA�Ɨ�Qh0���)Gj�{��eE����_��=��y����j�e���d�p�6�;� �  -J�,еT]O���'MS8#�����/,p-y*���#����;��������.kS��ڽ7��w��˔���X  AN��Û�9�f��	��
�)�h��)��{z�!����� <� ����W�}�9�=�I�A	������[np
 �'��&�O�;��;��\��'�+��c$���}	� ��Z��b�6Xa�M���!��@�^�KS�'S>ǅk�V����/�嫴Β�q �+~�ؐ��v����x+��9�Z���)�%O�'!�w�6�h�Z���s ����pK�'ô!�D���+�Sօ6�ib%��-��e�-�|���8-N<���� @@��`/^ %ׁ�&z�M8������;�_�`����C'�D��Sȹ�G����0G�����	D�M
�@�a�����5���xǍ�4i�;�8N�|x�� �%Ùw����j��O�^vdJ�q������'��&L���H�Ф�4���Y�}h�|@#0�4\�+�b�=M|P:�,EU��v�.���T��J�r���6��L-���W�Cg�qo�NU�e�Τ'P3pK�?�2Y��L��1����5}Q�������a�)x�
�x�J��\�C=4C#``�(�}/�v� ���<NBA^�O��z]���zPk��R:����'Y�7ρ�Ţ8�9V� �	�B�-غu;�[�Ě�����M�''�Z�R�zg�ȊP�N�ƿs�9���|��ch��#P)���׊�oJɕ�/OS��3L`�8@a�:��޲�z\�.�Hx1�����r�m����W�]��C{�O7P'�t��'������3&FNYɛ�((Ĭ���>���◿�\r~Om��}s)E�o� �<�N�1���+��Ga�
C#04o�(LռJ�^��8a�8��!y��*Ͻi���1]�B����Ć�ͨ��`/��^{<��J>�P�eeĢ�_��y��s�8[�������	bfN9���햮&>
o~/'�����=�R\4��L�!�#���=�F�Ў �CY@��`vi0�2�|������V�R^�J�
짟~��՛��lP������nG{�#���2诧����_lz-M��7m�|���Y:#'���	��g�2.wJ_�U2��Yy*�~
^�a<��y�����GB7Ѿz��eedV�e:t��������U+ �Y���8�����U�KE��_��f:,DzH'���Xu-�i�4�J#0o���������3�k��Ϩ>����4�]��h����O?�-�6��C���c��)�����z���D�NV�R2쯺�*+���?h�b� ����}R<f�7o�;5~��Z\�P����8�#0P���7
�*������pԘ��
ho߃��_���/�9�$4�c��4u
N�>�N�2X���F&�c��{v��;��U�b����>_|!�?���GG�.lټ+W,C���+״�]��/��a��=hj��_��r�.��S*��6"�<�<I�JA@:���;����Yu$�>��
)�W��C�d���f�J��ߦ����o����ys�	�T��=���d��*b|�ᇍ+I-���,���=�C�,V���z\'������L��p(�DW�v�1i�4�{�\�&�F���� 	#��b��f'����y�e�+��6K�[�p��cxk3�a/�#G�!ѵ;wnF"�i���c��{W'��rؾ'���0>Jb6V�_�B�yK���ok���3 i�#�7}�C�."c%3�xi�io�3�t:C��#vx�W���2�L��� ���q�����yZ���v�a�
;�>NN+z��n�_���N��X�a!��g�KN6�ö�q$ytv�p���4������� V?��R:iI^�7�������s�W�y    IDATq��{�����
�|�tn���s�I�6)������=�شq;
�0�m�c�)s���Et���R N�.R�ra0����[p�h��j����xQD��t�!���n�7�Շ���5+^��N�\�l\3��#ͺ��ץ�;*rO�Y�7��Q9���?���[:gW�<���3��uQ�X�"
�����](ॗס��	�mÉ�N�o�d�ܼu�%�l۲���{�J.�\sK�����m��o������!��z�أ�~���nj[���g�9�|7�n_�L*iڸ?@n�6�����6�cܸ�֞Q��_���)[L�z�[�b@O���"sz��E�����:(�;yq���(��\��o�i����5��`P6�ܲT����O>e��dOe"��(���iՋ?�$}TIHw�S�ߋ���ں6mZ��nrd�ΐD2��ϯB0P�ݻ��|���~�2|�E?��f�Y���D^E���������f{{���}�l�Q��cƖ��W��p�ٳ�Iw`���Hg%��:;��~�&�|�X�������C�`o�(jt��[]T�Ϲe���i���L���RJ�����������P(�����P=�`��hY�1N\<ܣl���6�ai��ʑ���I��fNl]��Mvu�����˟��܃N����jlܸ�{��J��o+WmD6�Ggg;v����/C�%�o��k�������#�Jc��1����4��R�N�~��p֜���Ѷq5�.͓����q�m؂L&�u�:p�)g�{��y���;��'�D3��6w����L�`�L��9*4Sw�����{���{��4������¡r���_��/��]~�=Nk�,����~���]�� ��><f��x|�]�4i4ZZ�a��W�˧��`c�4��+���Ua���5���n�����;�������imn���n�y����������-�i>��`dK3��<^� F�jB�Ѝ�{�!���y}~?��3ؾmv�N`��$\�vK�$�3��\4�.�"q���ӭC�9�	�����;	�n��~�LM>���c��^�(��}�ڱQ��.��7~�������;�q�W�ޥb���g�q����E�̚�`i�3`���]X��"�TPc�捌��G���;;�ص�\x	�=�D�bx��p�-�X:���+e�Z��/ۇk��<A6
a޼K,�3�Ma�m��ٻ{��B��k��<�gG�6lC8ڈ��q�;'��o�TOQ=|�k_3�gF�z2ݓ�AGaB���~`1 /{���6���A�zd�܇�y�ߐ� ,�_���"�̦3�\bꕀPU.��ty��M7�d�B�5l۲{vmEGG;�9�����l�p��֬݀t*�+���ǌ����nK!��������o�����?P�o��#�3a�x��w!	��&���������Ĉ������Z1�ē���	��g������ގ���:�������N�nQ{V������K�ސU���uoٹ����j@��U�C�痦"�h/Į��^'KJǊ�[)�bB��\����MT0���(�v��y������y}��N[��Z�I[Ԇ��[���?�2AҎ�W�H(��TO+D�5��i�0F���K�E(��3a
O�/�@L����;��{Cc�&6�{;�ʚ�R�����uEE�)�j�#�@֬�-���zy8��_����g�{S{ϻ�1��w�m��T\T��I��S3"V�~���<��/�͛6��/����ծ�u*�A8�$S̘q2�u����mہ��zK3�{�R����y��?���R�7��ۀs���ݍk��N\tх��E0�����F�����{�PX���b�'a��3W����R5YuG��6	]=��ԧ,��_�2��f�i�`ж��|Ŭ��������ڜ��`�^���q1�	U`L�`p�L��t}��4����м.c*e8H#���ܔ]t\3���@J B�,��+}O�ϟJ���Ϟ=��*�CA}�(K���^>�hx{[r��#�c����	�us��GY�p��[Q>��_i���t�h<ԉ�?���ΝkkQ���i}�ƍ��̵*^)i�<O���֐�U�\o-���i��IF6Ї�s�g��SO-�K՜j\U��yb�<��wT��~��`��E�G�/�������'5s�?���bʔ)`;L�'A�}�9�=ʣ�c�����D�f�j���{�j�
[�&p�>���KQ_7d#(|����Z��b��c�����h�hR6g)V�lʢ�'N�n�܈�H��,��0�� ��"",��Հs۶mX�x�i��(h+ �����җ�d������Y���H���j=��{��*Ս ��w�۞�@��'P��gg��-p<�
��g�8Â�
��$�%W��o��o6�2��o�G$�]w�mD�e��w�	�����a��s$�x�)���i�eG3��T�Y)ܴ|Ư��e롯���~̸��n�^��nu�i~>�����M���c�# w�R$�2��*�'����-�%�sK�X�I�����2��J�*�4Shm{�y9�V����&��@��~�T 4�R~x-u�b^�O<a>u�[i��`�`�x��kM��t�R�df�=�̳x��l���
�����[��_��_mdAr<�'��'L��"�t⬝R��'.f���/��K+�;�S(�����/�ws<�q}%�_Ҝ�C!ׄ��/���/�	<j�X+��ĤS�=��ng�Z�Ҹz�z�ro�>���M���}C��Y=�<�pT��i��]o��4�ú���4<��;��P�������*�Z
L��XȦM���8�K����c��/8.�P�|�[߲":�6��κ�����y��n���sx��|�,
�����YL,ܡ�ƹ�Vʟ�'���P�'����:Ӧ5!W�c�����'>�ѣ� ݝt�鴍g>Wj���~�,zx12� ��"��&���4�\c}��$׮_��~�����3�
	�a�?�S����Ϳ��q�1��nPo�y_뀱�5ZT�����߼�M�b�}T����*;�DkF��K�Fp_�z��w�'�t*z,� `��:�ݏϨ����;�-�<y2����@��2�@��d&��h���x�������y���*��d�m�w���?�wį���<�M��/���b	���aĈQ&�#W��c�m�b�H\\�r���2k�,�`����	&4��{���{����a ���X��k��|j!��%���9K}-��	[�)]e%u��i����oV��y�j�/^���{���J_ڧ�Ҕ)|9����%
�4�e�!����q�Hx	�5��X 3�.����b4�K^��||^��8j��}w/��9�т��z;Ə��ꪘi�Ŝ�1A�߬�l��N��~�%K���b96����80퐂����y]�?߉���_X�̲�<<_��֯\�\���ϟ���>�ƕ��j>��y���J»�:��B�2d8��I(��k�YY@�5 k�d�RYܡ��^UV�u׾����rl���%v����*� ���SӦ��jL�:3N�i����Z�\�(�
ؽ{�Y�_|˖/�`�Yxp��IH�ߧX,f�[Zo���^6�����W�` l����h;%-?2���}���b�č� 087�|y\�
Ԋ�� C�+]�r��Փ��:s�L+�b�@n-�}�C=4K���"?�Lpj`|~� ��ǟ\���h�`z%�g������ K��UV�5k
��AG�$�;��I��97��xg�mJ����^ם�W�����1�t������T\O�J��}!�PЇ�G�D,Ze׬��3��s���Z�w2�l=���� 	���"1#���lr����u(5>r7�
'6$Rq��Fg/�*�D����1�y�ǖ ���WZyA��N��8����\^|^^��*/[��x���Z��ť�����.Ɯ9s��X������~r�0�DE���U# ˓���pMM-fgry
��)���q�;�]��/ 
�?�p�T_�Kk�����{��_d�h���v6n�w��:l��6`�~̂�a�	|4u��5�F޹���h\,��c0�~UnP��e��dpL����IVgi[�78d�3���M��Lݔ����H3���+�?e-�R��@����~�^KMA`>���	�y�,+l���u��y׊e����r!�{�����5�.���u�}|��<�"Zʱs�Nz|���[��Cw:�T&mY�W�;m��#����!!dq-�)�l�("UQ*~'A�FD;�#���Z�^7��-ŀ�:Ї�?݈��y��'��\^��)6����-�,^�1�Ә�8a�Cʅ�C9�P�"�����82�ɖ�,�8]|ʝ����&L�0wkIY�4�C�_I�/2G��l	���}6�����28_A �w� ~�}9�o�<��XNjE�C�'5f|����P������O��@��p}/_����ƔF#w��@��m�k�C��8�jb�ո�	�x/�W���'���=�Q�,�L��|yms[T����+뽏6�4P��xm���_
Z(���x�Q�o?y}9㓊R������w3Ѐ�(|�XЕL"�ݍ��%BB>�57|F>��G�{��=��Wf�U��?�nP�}Ya��������;�0J���T�Lk��O�TP_{�{}	cY\����|?zo)�^+���|q�r��w���|���:�ڰ���,Θ���w�Wpk���ܰ�C�8>-�XUM)�9�B�Y���ks�u����@n��>���Uޏ_q%߾>��O����j>.�o~�.�\^��b�t�wmmm��HM�	�|z�q�ۥ�b����w>������c�F���8&qӊ�n|����&PB�2���9����
��	��1�j�����	_�ц�������]6P_�� �E#`?	�;ݎ��,A�� ��է2�}��V�[��|pL-1@<��2�4~���ZEWy�5�׼{�Mq�}
��ރ�Y�W�e-����y���t��Zpoփ�8�R�O��SƞR_��y�A���[0�g�xǵ�|�}�������k�k���11��c��w �G�r��R��w����'�&��f���iԇ�k���m����*ȕ4z�p��#����������Q;��W�ل�G �{�B	�$ zP��i7�_6�����{+��9���WC�����aN��{�B���L!fŰBPy��'�Ng|mK�������b�U��S�0���@�����;�C��k����iT����*��c=އ!Ϳ�ٚ�`�/�����^�/W�4x�b�?X
ZQ�C�!�]�J���K�0y}d�݆����}�f=�s�ұ\��E2�EE��"X6Iݜ���S^�}	�y]� �==ǻ�D>�5��o<�~Me��_�����p�L���h{�Y���8��K�;�w�Cm^��R�@~�ײ��!�?����>N���t���b)�3�C� ���>�`	&�B5����|�S!69���A�?�~_�P�˗�*X�0�$ �R�	�S�2�5��e_4����!�?|��/*��}z�?��l���3�K�O#������p.������e�x����W
��J@����A��3o@Ϳ�p9��.�n�G� C����uL_i}"�� P���ؕ�/����^�UX�C����:ʜ�ޚ����3��f���r�i�o�n9�{[O<z>����{�!�<���_(��1��7����qzh�;I�$	 �M)�._7d.Vs*7��+����a��}\@]�CK����+�?}��Z:�?h�>ݩ��;P�t�!�?p�}�a½�z����U1�� ��-����[���om��`��-X���x��*���A��9_�:���W1o��0&�������h
�L.�M��������G#~�@��+Ư"Q7�U���U,���7j(e�0E���������"P�~��������ZB���R�?��q�|t�Z<��*�Qі\i,2�Y6W��Ze����y.�->�ݔ���1�G�����0�^�z-C�S E�9s�(�O�U9����nx�p�d7�錍m&�~P	QV�����|V�6���J�9Q"��p��*k��s<ʬ��b�bU^
�ǎ���X�� �k<�TZSz{+�5��ޞ���Y�益=�{C�Z�'�jo�^Q���G�\�-aV\>_N�渲��\=~ �h����=v�+N̻b�e˞7�qWp6��?��y�"���������q�?W��E.m?F�����zm���>V�=�B!���&-�j`�&K��k�8��*�i���#��?��% T0t8��\�L	�ci���w������n,��R+T��Whv�L�6���U9����K'皙x+O�!is�oW8�tm`iS(�"/���=^��J�������E�+$^���������r�����@��)巪^�hir�Q�H��.9��8q���lh̩�X�TI��
�%�����sz]���~����|g��8�t�QPp���sq�xoS�I��kk]��������)o�s/�'��Ϥ�=�i�ڐ��U��.\GV�۝Fsc�1�2|ذ$Sd�u䆉�k��V�$�[���9\�\M<�p���/��m,G�Jt9���g�y.�{>��r�O:�4nFiuiv_�۷�4C
m i*� "��F!�	���w/�x�B�`��F"�i�RW�~��/�1I�Tۻ��	��	V��x��}P���N�J�7 ���#F�w��W��ss.�R)mb�8���;����x
x�Yc-�d667�S��ל���_ȣ:Ve�.���pu �Q4��
"�c���Y.���������:3-��E�,&	6�#��(���	N	X�{�ݏs�{h�Er�k�;����Ha�߇�E��,-	j��Ƿ��ގ�=^
/��'��s%���g���0�Z���ӊ>aډ�����W�.�h4�ؾ�:s���T�zV�X���q�Q��-�@�ɞ���/����x��>�>$v�3kcU��e�I3��oKS#2���X��Yk�F�-.��ԩS1i���k���.l�B�a.|.n�#�<�ƍ3ӍVB���M$-�C�?�:��~ ��MWGg���h��_<�V�	ۻ����{r3�1������ �U�oV��m�L1	g��ZB��TE@o�W�KSK�Ϳ�CZ��xe�\�Qy���w|G�]���Z���ޝ�_Ȥ��҄=#���]���=w����!��RG����f-!���Xr\ml
���:+a*ˇ���J�)	yZd^b;���8n|w�I�=	��LyǕ�	]�	bY�K�P�{o�Y�)���:֫��~N�:�����~�s����r��9%(�F���q�U{đ�DB�fRض};�y�i�w��Z�Ţ��;|�H{�h�Ŀ�?��'k�h�i n�A����a<�qc�oմ����q��ދ�G����(���c�`˖Mf��������Gy��v2b���nH�L�~�7qQ���<�_c�@n"i�2����5�v�����˟1o�E��H���|�I<��2[%��ߩu^xᅶ���
8R+	@���&�Q�)���x��)�i���8q�]OZ�W�P�}�=�II���^b.�#�l�C�^j���e��r�xP�����;y�P��B-͍��c�8��+7倾�]1�<y�]w݅�/�����F&H��ƙk��#8_����[��yK_x�>�h��D+�q�e��36GlIK^S�7ޗ�p�w�y�)Di�_��O9���J4^��uE�C6���l�Ə,$�}8FrG��ټEc��,Y�[n��L�,�X<F���1a�8�
i��	,~)^Y���&0�!\g��L���3g[G&<��_����j��F^\�7�s���?h��?�'�S�.����w酸���+f�N%�f��xa��,(GL�O-lW{J��s    IDAT��������r�����F�L'����6�}�Y�[��� �!7�c�=f���J�����;�k{�K�5Ea�9�6��K�$���{���\m�����5�\c��X�x�cC3�{��6m�\�*�F�v+-��8y�d�i�r+�Y�.
�qd�1���K�N�/�7�bw,cW,���s����c�<�쬪��N���IH!	%4�]P��2"��"
D�*���S��\D)6H �t, ��i�L&m2s��~������̙3%���'�̜����~������Q���ި a��}6��{�=���FΪ�j�p�~����4Z>��#�;�����f���Bs�8���2^��/Y�T[.ug��Y�|G�\g�64���˵��|3~uS��ڧ��ֲ�Ro��#���4S�Y����9R��q{)��T�E<�|����i�(Bt�y;J��J>�!y�'���u��qo(�\p��Cy�S��?����V��{
��"�3�.���mr��G��%y��X��t��Z	8���e$��� �l�Pe�w�o&��^q��2k��2]��c�� i@���Δ��6Y�r��tw���<��w&,�ΐ�9�<6��p�X�[@�Əf��~�i�%Lb����!|m�r�є�i�����y�W�blsr���qPbl�{u_ɺ1��5`��f7���D�E	��ۢ+��h�ԼV��i��9�����g��5��� �W~�����C�h۠F{�6|(���i9h� �O`�`lX�?��������t���K/��ӧ�����k�W� *��oֱ�/���	L���s�Ygi�l���1�e�*T��9��́�N�lNۏ�X9�kZ��0��DkHU���|�u�i���|��k�T�� �Fu۫~�k�g�ش{�=���|E׽�]�y��=~?��hw{>�=~�}③ll^,�T�������˜#�X�(/��5M�$���u媫>&3g�.�lA�x�or�=�H,��}n};#]��~[2��J�j�O�� ���ڨ�}�r�����r�rI��f-�M�NGd��9��cK}h�������	�S����Р��CM��S���3��r�����8E��̵r���1c�>����#o�q��hO �i{h~F�������K��u�P7���q�  |��6W�k��J1�b�?�^54f�Q������yJ4E��q��&(��Z�v���_j�E����瞳w�/�P��t����E8��Tł������ G�q^�*��;�MPs ���35�ߴ}s�+�Qp�6��)SJ��	_w�y�j��h��Dw���t6�6׀?=|�^0��7ø�m��+��_���9��W���UysچR���i���ӟ�eie�yN�w��Hn�g�zHƍ�˸	�d����U��tN�-]-�\X:�S�����sϒQc��ˋ^����_��͙;��ɶ�+�?�3,�ٻ�&W_�!���ic�<���r�GK>�%MkWIgW�ĢԨ��斤4�k�l6&���d���Ҳ����җ���'�E�hٴ,$۴��'NP�0-�4EӺ�Kܞ��s����cƨ�vb �wM�t�E��pԨ�ȖIH�ײV���h�f�"�\ )���`416\_Z�?�/�B�'�d=�����E��s~��|l�an�]��/��8-LШjh �1�t���CF��o�k��8�]��q2f�o�ͥY<G��9}���ic�o��8KN�~�X���J�w��-��x�W��u{��W��c���uO�ߡ�� ;��{��gk羦&GU�u��O|B��|�+�'#���3F�,}��ڰ'��c����"�iiMI,Q/����$D�I.�ma0{��l���G��?g��&����G��s���#WX"�����By�O�!��-�XA֬]�m1�
��l��.�6�O�F^^�V=�(�B�(,P8bQ$��pL�����Xx�Y4A5����4__s5A��-n�O7��1�	Rv^�����67	b�e���>��kn}�ôG]��xWz�:��1���� b�c�����>����S>���'��ρ%,q�\�:��U>��/�?��aB����� >���O�z�{3Kz{��Ӭu��>�\N#�h�������{�.8}�~��l}A�]q�J�-_��<��{�G�'Ə����)Ţ�ĥ�+/˗5)�l��)�Z;��o�Pԅ��䎟Ȋe�J}�s[�����j�Oz5u�NS��k>.�b^��.��m��c�L�]6nZ+�=�.����d�4��$�y�ؒ��{�E���*~4>�i4`�J�^8M8P�p���;��1���Ȩ��6y{.�j�f��Z�@�`*�8L�y��}��7�EE��iަ���>3���=�����;����Aɿ�	=�,�����ܒ���(�&����k�v.��]���+ 6���o�3��M �
�	�Jc���߿��*�����s�������2����� ������Ϗh(�2���X�PfX(��׭�'{P޲�,i�8ZV�y]2� ?#��lFd�+�K$Z/�YIeC��]'��Uo��fY�b����R�Ap�������i��}��1r��?*�u52nL�,��Sy�>�J����u���ۥ�G�	i� �[��+#k�&��S標�Åޙ?~ɁH��SN9E��Ǎ�R��[nѰP��\t�F[����j��&f,o4�������L0��i���f��`?_�5'���K�F<�}4��9���h����(�Uic��H����l�|6�v�6�c�='��} �4�V�Uc��߿����)��l��������}'�/��y�fY�M���j�f�� ����9��w,,z_��X|��ΎM��ӏ�N�GI"�ի_�Tڕ�A{OO^^|a�D�d���r�ۏ�y��֤?��w/���������3�gvĂ�i�7~��-yU%ڇ�Y��Qrּyr�[����VI&7�����"�0 �➡~��Y׼Q�6o�T:$W|�*}`<�[o�U����׿��=1�h�\r���%�m���.�C��k	_��,zc�x8�/�\��4/_����/[���[>0�Z5�� ��7 �/��|喏��]������<>�җUe��K8�}k������J��ӷ<�}_Y�����6��/��p�z��Z�׵G~��7_�~"��?�|����͊�Ә��@���j����ѾQ2�N��R��C�����BL򹰼��5iK���^";�<SCA~�a���%��T��w��u�=w�}{����/���xC�=ye%�ϓ��T�n��v�X$������MR�Nm���K!�x�N�;�p�m�=�D7�勉ǂ��K������w����%���A9j��x㍚d�S_���y0���Q9�].��V3�r-��r@,�0 ���%`/&tʩ!Ӽ����W�����������2��}��\�3��e�F9��[ff��c����W����TK4�ݗou���r_�9�4}�����$`����Ja��l��K�'���p?����K.��2I��*���חȚ����t9k�#TN$��ttfd�Y��A���@$:.��^eFՎ���77�a�e��Ͽmā�$/�_#k�9�t֙g�	�'�I��Eem�Jy��G�E�4��E���C<DN8�d�0q���&����s>��'1���Q��	���-Ġ_w�u�v]�j˖-�gc��e��+4��6������26g_Ԑi���� �\s���G����1����s�F]�w}�5|����[�3��)��@����?._A(�r��`�mǚ 1N��90������1�[}��h?b�W ����XC�w�;\ߊ��Ӭs�s���WK�K�dlD�� ��<���}�{�+�|��c��j��_�����4�]��� ��g��M�9��s�}$�/j��G{T��կt�`�/pM����M��p����dā�����f���*���k�/��޲�d�i�0�����.kׯ�H$�^���Q�'���x�F�v{�-�76 ��,��,:�a4��{�q�>,6?m~��w�߷LO�2��6�m�j������V�7ЄmL�¡ڵ�|>�����7�-_p�S��P�Y۹lN�D2~8����1�9-⬿5�h�Z���i���ߟ�r���{���)�}�A���5���kв����w��cʬL���a��E5���:���.3w�x$*�|J�I(]�\-�J��<C����Db���勲x�k��L:���Ek)���;�~������)h	�?$17gyW���c�	z�n3R,��ڶ�X��H\6lؤ�(�`8{��q�<c
�>?1�"�.]*].�Ӿc��@o8����w�\����\��U��>ܱ�����w���	Z��\)�u[i>�\>������KHM8p.~�4q��}�9��{Hm]��pF�Ơ�s���W���ߟ����w�a�}/����
`���T؍	r�TzB�ϸ����d�ӴD ��<$.��W˚5k4-�� �Gc8�st!|�ߔw��r�W��C�_��7!�?����0��l���\~��-^~�9c��(�.�n�3���1��3P�ӱX |ƌ�g�$.�x�����߯`mt��[��:;z�V>��#d֮��J��m<�%�)����/��ؼ~�
����:�{�
��Xο��kRa�]c�b�uM@��3g�t��ٔ
2��E ��n�KI7��'�"c��D�|�T���p��iZ������V��b|4���YMPq�JiB���m5���1�n3`����ӸSj�S����Z�T�%�+�}OUU�^@�6|��h9�F���)Sd�3�&Ӓdv�x}�J� l�����ߜ���\�ol�)ٞ��R��{(��n�� ЇM���+�f�?U+�j�HfK�e�=��h��=���t ,�`���{�Z��~D~��ȢE�Jac`���l�d5�,�6����T���lc�{ ��ߎ�7��~f�PoW"���ֱ�O=�TU��A�ɜ��`��?�h��|�8w-��)���}��8��	ܾS�x9��jUϑ��6sa.�9����s�Ľ{ci�����a��s�2~��7��Q>�yv�Z�.b�����'�"ف<d���z�qu���ʬs��E�7i\���6�q��ގ�w�j��MX0C���Z�r������O�'�?��u3�9W�y�1\3 ^vL$���G��� ���w�+�F��?w���d���4<��SIO�>�$�o�]X[X ��kSP���9UM�дa���Z�2�V��pJ>x�AB"Na�},���!}����i�&��~�-.,�-��������������3��g_X2�%l�!��\����J)=y���{���U�H6�@�I8fmb�*KmM�*\q�Ǚ�^��M;�#B��#����xK�=yI%��|>� O{�z�Eh◭T��{�("�|o-u����� ��_ViM���a�QŐ���'�/�o�m�X��p��%�X}|?���E2X�J���p���;f��},`¢x�ꯖ=nܻM��('����5�q���Vp>�f:�v�D��������Wp/��\��B���,��3�4�������8�*�O�n,��F D� ~H�0���F�
���j�Y�u�c��'�.�����c�@����]�\��Ec��p7����#�4ݓ�s�Q?�EE(p,��M��Ꭳ��{�՜&D���1#��}y�m��a�zO)ʡ �bX����tc�z<7֓����	u��w���T�����g�r%,"N�{�iڼ i��^�Z�
7
��7�Is��G��d�?tE���\�4��
��.�;�R��Pi&�����c
"L�N2 ⺨9M\�GhX�
 ^V����
)dz%�����m�2�/+�ZB�{�k����Z�6���4�+>t����Pi)���L^���9��SUU_4�5Kry�21*E���D����x4��H��Hb���9��3���MH�<�Ũz���ϲ��֞�H��	�hB�Ǣa����ϥ�~�K졭g��o�˜�VEV�� yʀ�֥�_�)��o���xn�G�>2���
Ղ2S�d�}��P>4��!3�%�0.	���}O�\�v��sP�G6�W��#!��b��$1�,�6��� �Y�]X�E��D
���F�����-��s���?f�I'�K�w�y������ӱ�5	m��|J��X �>������n2�`&��8Z2y���$�1	�3�tHM�[:�֋d���HݨIR��%��c"9"������ϰ�Q	SS�%ߛ���l�N
Q�LT�y�Q+�ܲ^6nZ��^5-�C���~��d�`��VdN�.�ϱ+�3�����7!�X,��>��-�ʔ9W&ȸ�j���;����p��l�Y��`���9����0]��J�*�|���?�aҥ#��Ϗڒ��*i�L:@��C����a�e2���������g6�.Y�����r��6�Z�v�g�;K�O+8�
y��@�i��o���f��_��u����/
�c)�$ �m� u6��SN9I�<{���Qb##�IL2�uHw�
y��dݚ5���mǾSƌ�(�bA�E<�0�XC �<�
��Diբt��k$'��8I�k$��H1&ɶ6y�OԒ݉�:�Td���/p��̙��YT�$�Ȣ�,�k����O�����DùJ��	'����{�Z.e�s�b��}�����e>=��h��M(���zA�%��{4H�T+.PB��2A����_-��'~�i���k�FMM�F�(؇c[4Y/E�� �B�F���˼���n���P�M�I�Nш��e`<�̢��;��=)��Iy��h�#l��\;�l��Xb���!���*�l��J�G
R�I$�*��:���Ț�Kd����ݍg�����y���6�m��d�*Z�)���J6:^�?C�z���i�I�������vB��'�r�c�� @ȳ:�3�$	�>t�	&@��}[so���$f�(�ǀ�$
�q��aaS�B��������؀0N^��P= /�5��C�R?fQ���2�SJ�?��[]�o�4��YҹZUOʹ�)�ȡ���ۅ[9n������b��L������+�V�i�,Q*%�˨��F]�Z ��S)�ɤU��L�H���t���-5��&"�#t(
Ю	����{�±Z܊��D� �\���I"�"�^p�lްF� O>�Q����G�F���ry=����c�}$"�P��#�$/����-H}�hy�EjE�ui�x�s��{�� {Y�y��2�47'�>3���g�f ��Y�Ͼ�i�n��O"��XY��7�կ�ϱ��@ྍRV��r�Vp�ņr��ou����J#	8��ܵ���c����;��dۇ*�>,>�4��:�ҮA3�#�6���w�}4������
h"h&hZ<L4��1���M|���|�v��U���%�؈�	G$_�jr�Y/�x��82���wu���qN`C�`��c�f=|�J���*d�.���P��:W�}w�"��keڔ�2g��R;a���Tt�`�/�׹�)�~V�DX#��IE�J66Vr����b�F��H��I:�s�x�|U��P�7��8�h�Dv�\Y�4�ӟ������cL�5���&�:�,�����k������?�W�u8���-�����d���RS�ڻ����h�
���~�D\B&�SkE��׈�j�����N4�|XT�pL::�d��3��w��͘Q���1Rp��ާ�|w�,>�i4�%����Oߏ@���Q*��%w�_�K,'s&eD�D��gs8<��Y%C;@�0�H���p����3��)��&��i�f;%�k�����n���52i�$y׻eB�N��I�)��I<�W�@�O\�֑��|1,�P\ґ1��-    IDAT����Lx�d���
jRc��7|O��Z�B��r,�2��G{Qd2
 &<�֦�����G}���e�����G�{${�,n��u�ܹ��'��)K�B�ׯ�iJ�P�����Q=%� ��!��|��r�1����SU1����ē�* ��]J��T{�#��5p'�V�,׏�M���#o{�12��4M��f{4�C��_A('��P(��1��'�����vg��o�|���a����z��|Njh�I�i��pF�|�'`�!�i$'E�hS�lЧ ��n����@ ����,�^�7~�g��F!-�BJŤHO��������2m�t9餹�0e�tt[xja����POH�BB��h�9�	�M�j$����z�>C�߰a��薛�E/�0@�V�۞ c9! �瞫�}ӊx�-&h�ϛ��|� (�ƽX3h
�)��Q�*f{=#��L�(:m��ɹ眧U=�����&�F՗rn ����0�A::����ğ�T����j�/��dD�>��������G+�>x���h������|@b���]'==���+�i�Ji�h�D̳=��Kf�ds$m�f�7�t�.V���o}?���4����[5I�c~=�<��-�J��R���-?Q�?����Ȼ�}ݜ ~�����$���4�����w{�?��X]7��#��vi�u-ᨙ.��%^h�pz�ܿ��Ҳ�I�N�*'�|�����d�]D$L@��7�gP?�����? �/D%��tt�d��[/�P�&|��ٞ��������R�\���@��̔+��s���a�DЖO9�Ufx�[���<s�G��5i�ja�>�VC������k�[	��4t:pN�x��ަ�N3���e���I��J(pN�)@�˚�����YH�ͭ��ZP���=r,����#{��C-r�N�;Zeٲ%���0y��m�=eԘ��Jgg(�L��ؔG�Z.�F4��il�v�=��J����l&/ӧN���u���mw3v��\�T^~�yy�����E�A�%@gƴ�e�}���;Z(���z��'���]�t��g��P<���L^� <m��kl����a��5�7Ż��U	�K����$�RISP�����XM��p��%W�v���I1�)5�#��&��*���Ҳa�����O��:�cͻ0ϡ�4r)� ��>�� Ӝ�I&2�9|#��KǶX,!=]���?��!I�9�a8�>>�E��U�X8"d�J$�O���0��#�=��$�
eb˾cc亥���w;�ʐ�&K�4(,�p�PO4� }�#?��?��pn���_�Ĭ{�@Y�2������n�:�h��y���?��J;�C5�1�M��e��瞑�uM�A��tugd�]f�G-�춇��.��GV�m���9��w�?����B#jf��lZ
��,ym���ҳR(f�.�~�$�HWGJ:;3�����G��
��w��]u�(؄���g��?��j.<0u�i������g�yF��玚��x���P���L$H�l������m������s��(��P�S��Pf���[�e�j����j�)�?�揀��Z�B��֬Dk�P�JN�%������	��p�v�wȝ?��<�ğ�TW����۠% ����I�����wb�)*� D��c�t_����+Y`
ʶ�~�������������}�$Q��c��|���dJA�B�/0�J1�W'k&S����䢋��C�=�~g�)�����ַt�~tc����_�4l�����^��^]$�m%�^'��:I�����#�~�z��݋P��]?W_ k����0i�#2�s��9�J&�?^I�g�y_{����.�fH,"����"�F'��e��l^/==��$��rE�ܒ��%3r��)S�(x[M��i
\�f�Gu�nD��X��K��అl�}�-��K�`J����$�$ �A�
��)���}
P��JZl/��UMG���4v��%����������e'h�������0��|�o!\�"Ų$_�s�ђz�6qٸ~��z�O��?�4�m��e c`n`=����k����g�r�Ъ�<+V�(Պ1+´c�?h�"4��-4gֿi�f���l��QF	��Ϛ5���D׻��V>�����Y�k�>X����(c�D0�P�$��{�{�k_�����8���.�HA���p��4��/�X9�I�tHrs���6˺uM
�(A�C�>���^�^:���K�a�Nz����k�#�}�'ߑ�z���%���l~^�N����5��6�{���v���e��W��#��_$��u�7K�ڍR��,[�^�9��ڸ�M�"�����d�����f8���|�C�/}�K��iM)k�q�8���CY��!��d���z-E��8οv��
��2�k���u�����餝�{�	�L;%Z�,��*���M��NS�?N�'c'L�t7��f���߬\��a�0GaM��b.�%%��d���ʈD��i���G?�%˖J��m�/�P�`�_�������X)�A�Y_����΍ՊF9m�4}ˀj��9�ǚ��?������6 h��Y066�T�S&�	]�N�6V�p^&P̪�s��u�]'+�-�4�cY��%���|�;
�P@|n>����o!-}��2u�x�PN^}�F���¡���s��2v�N�t�j9�'ɻO��x�Ң�jo�,ݻ��_O;���/�s3��,���c"��l��$���r���b�G6�4K{{��c%.�iY�n��sY��]v�uO�n?��M��/|��ݢ�������8�8|>�я
-�xX��o�߰�]�~�W<�ޠ������Z �_5�=�/�w����U6KK���c]���'�3�����e�r�#�|U�'��������t�<3q��)��eu��3;Dy��D]M]��Ʉj�G�K6<J2E���g�f�*��?��Mͮ�S�(7��_�y}[�?y&֏��8��;�	 �~XVn[�&\��� 5����8�aj~��9�� ��bV�YF��=7� �?zf��뚀5*�_��<��g�^��Nj,z�(=�Qj�~�U�Ę�@��n^/O>z���,;�N���AW�?&ٌ��Eˤ�v�4��$u���ǯ�V��FIgw�^kŊ�zn~�����h�l�0�k���CW^!�pQV�\*?�k9��äP��VKWW�s��jd��ViZ�IB�zY�z���!�)g&�5�\SZ�,z{8ַ�
��ޟ$R��8�m�9}�`���s>��� V����5�	p�u���o��匇�EI��֑���
:�!
B-f$�k�Da��3����&�}��ɪ�O�?$!AcZ�?�H�\J���7,�bL���;!���_�1 v��%Z�aS[�UE%t����mƀ&b/Ӝ�Й��|�R�P�7��zt������$8z˜�s����\�	�q� �����H;�()s��}[�:�F�"�L�.9�i�t��gȧ>�)u�ҫ��k�U`��K�B��&�h�x��e��k/���J�<r_i�4V����1���l떥˚%-׷KgwV��m�caٴ�EE�.ݲ_���Vf�h(4�=gϖ�\}�Ĵ�C�����;�y���]�~�jimkQ隈�K��NY�z��r1y}M��e߃T�ǼE�n�Q�>X��ӊS���Ik(���g	/��@7�v�cK�qmAT?����\2W��?�}�� JNi����^�+ڡC�������?�q�u��LN<��D�K������|�.��?~��h4RD"�!j�Nϗ��d%$4 ������}����#	��(1��|G�l��5Do�������M��F� �ti@���}�!��1^>?�uW~,�e�o�I����_�m��˵�"0G��6?�o%�IO��í�i�Ҵ}_0r?8|���<��#�<R-�;�C�.]�S��g�(�����<����̖q�G�kK��K��D��saye�r���ٕ�L6,���:=j�tv���C��0&?:�����n���5�5������~L�j*f����ˡ�'�b��Z�B
���i��M����뫤�#/k��ȱǟ��?���8�j4R1G�q�<,6+&�]w�UJ��}����M��^��m?k:R�R�4.��k`rSBAk�����x�C��崺'��2�
�E��ˠ����Z��K��#WKD���f%�k�p�E��M�o��u�d��i��O��JW� ��GjS�;res���Y<9��\l���%-=��C5�'��W_����/k}�����WU��d���b�ͱ�),�}_\������[Pۦ���%
ڒ�ݞ/�K@���S��,��^������Fa��^��P�,��PV���8� �gs�Z����(k��a��iz]:�h�p8"�]=�|�jIeD6o�:\�8���+�_[.w-�/�5�m6���ܹ��L�]]���]�F�{�{������ukVJwOR�6��\�Gyr�$ź��U�o��Y���רs�ŀ���4v��v�J�{�WZ���A{D`��㎅R��s\s�j�O;.��JN Zd,���u�>���xc�����Ւ��q�:)3D�E���u�jA�l6%�t�$�Ih�g�Hj�<xϝҺa�L�� '��Q�O�.�T�GE����{�i���	z5��aL.2Z
�1Z�!-5"�z�<����_��������C���F�;��sh���r���A�<���a�>5����l�}��6����oK>M��K��l�K֭}U2=mZͶe�&���n�hm]��^�$[���ʵr��W�����p�N~��?�/�KF�%����m��8���m��+���ƙTJ�._���$P��d媥�|��QL*,�t��5������3%��V�1swV$?mq�qN�iF�C��x�%n�E�B�s˜J��ETqkT a�泙��:���db�5;1W�=�5�kj��'%�Z7��U��?�u~��-k��1�[�y��w ���F�eR��vK,��!�l����r��ۥ�y�4L/���4��O��H������<���2�4²q�a)(��B�^r�1*z
1	'F�g�)��w�-���Ev�?�����/�}i��Q@��?��X8u�@���9�9���/��ژ�3�����M��A	%�GK8�q���7ȸ���N)Ƥ�'#>�;��?�s��~��ɫJUϠ�b>���cG�YgΓ�;X�]�m��i���7JG[Ri�P!$�h\�L�*���Qv�6K+C"�)��׿�����x8�}48U� � ���4�����kU��*�O��q����Z0*��%�i�OKWG�߸�E����$	�Õd#;���@�/���S��f.��{�w��х|F����%%�L����_�*�Vj�ƹ�d���E���lZ�ZVZ�IT{���/��/���I12Jr�Z�)F%�-�L^�Q��ǷH"�V�v���b���,D��2F��GI�)�����w�h�믿^�=`N��7�B&5��x,,�L�<��S���OHw��E�g����Ւ��s̱�����3V��^�Q_KJ���������++i�tɱH���0I�s�<y�[���DL��Z6o�H��+V�����HmM��7^r���?�L���ø@�RY$h�˖-�Tp�r%j��vq왃W��ΰ��_� s�r��O>Y#���:"�Y�+�fZ|�UWT�z�5�O�1��<�v8���N�����*g�{��I!��P!-�ѼD�ݒ�l��~�lni��;M���q�$�FK���Dj���ϕF8�5��/Z<>�0��:)D�$NH�>��:���R����)��H��ڧ�2�w��ه~�nԜ�D�QR�`�|nV?�d��Ib�߽�ҋe��	l5��sҶy�,Z���\�R�'64(1z�X]�������=��qB>��_��?w����+*�?tN	�pxf���w�q���{�)��u����%� �ߵ�u��IgSZm�����-�>Rn-��+��� "p�P��/�+�A����í����ꩧ
U�Jt�g�����|�s��д,�?��I�=�y}���~*�%�&M��ft�m⡜�r)I�Ҳ�y�!p���S����K��ه��O5h��<��#T �HB��I���ȑmIm�M�em�j O���Ù�ߡ�7[o{p��c>9����M�+�y����^�����l��o�8�!� ��sl6�ў�T�em�_9.��+��������Sa��1�uw�q����46ޔlO^^	���IM����Ak�\CC�w�}�|��%��C(�鲓��K�_��,~���q�\�߉r �k�]w������H j��3����@�[4�j�A�ᆪq.�K��h��VD�B�}�1b���E�S�`�M�X9�� �j�ѨjN�\A{&S<-��Z^
�n���G�R[C7��� U"q���?Q���$��Ȃ���91�XH�X����G&�W�N)�"�R	�X�n��/�},J�֩	�сo��/L @�@����~s}�].��6N�i�2(��f�TAA�US����fy������N�����r��i���8����HX,��.$+���̓�8q��;Fv�4YƎ'�LQZ[��ҲY6on��x��f|FA�h���O>���illT��駟Bİ
 ( �~�����G/m`n�DS����@�NA��k]i�����s�nL���D#��N1��
��pQ��٣ɴh���ҔF����fc�*�e�xI�Y�G4Ɯ>�Ez�F�bk4^��c��3��(��ZKH��[�C��ܕs{i���\@ohhJ5`�*{��k�.�{([w�y���`_�P�~�����t�"�&V�J�n���"��YY�v��X�\�֮�J���Je8�S.���z'�[�gNc�-���%�4�^�ؚ��"�J@K@� +@`��"���ʩZh��l~��Ԇ�BVl�c�.���`IahF�{ktMY7��(����B���-�6���)�ઍ��E1��r���"EpÚ�[Q���h������x�P�P@e!����I|ύ��U*a�`�--����`q�V��O������'�Y��	|�����Lk-�vMS��������5�<[�4i?1��k�߯Y�ܧi�(Y�� ��Z�~�i����I�$w���to�M��?�>�����̿u]3!���YG+\�a���^T_#�g����Ȏ�N^CE��j�P��ҕ9��<@��tJ�o���n&Ο�Ë��;�s4������Jv��	zr�i�Gi����F� ��Z>����| �WH��m���!� %�+p/}��n��p^.z� 	������%V/ޢN|�|�1XL��s~9 ��FeP�pŅ ���=h$��mnݢ"��Kz,�B.�^B΄{�롅㿢�N�����˪�Z9
n5���z�)���u����_�@m�@f��,q�G�PG�:��h�֢p�X������2��:��]�����ޖ�����ی�i��)�
�1���p1@ӌ� �@���O'Q?<|8?٢p�֤�<�[h^��]��Uz ���瀻W�@_-�-^[&ܠǀ+��ZVV��IT�e-�$z_N������c����7��'�O�:a}�R��i���[-״{��
h�\ֵ�t����,b�Y��+_<�ׅ�|���z_`��û���,�J�P[�(W��qƫ 3kz��a1�~��&J�T�=|���A�?�A9�c��K/U@�o�x8A��"G�h�Czq��r0ƔI���}�`D��@i5�Kt�o�M;���(�JZ�3�\sj��X�l(8@�l67�  O��
�ق��P�[]4�7��0���5|[ݴ�ܒ�\��`ӻ�x	���m�KTSp�����?98�X7Dy����~&����5��E�JQ;[�oL)��>��iHBt�����n��Ÿ�H�p��j���:�4�H    IDAT^6�����2�+�5�K�'9�zDd��b��c�ҺY��j�X�{3��"�'d᳧���Ju�Z}.:���#��t�9x�G��6�6Wt��+; ��`�=[�}|�|;��_�K���7.��V`����n'��3Yՙ��d����fZ�{u�Z��>ڲU[��>�?X�zەuc�����7x'h���m�WI�!ʧwc��p��1�w[��J���T^Vc��%�k��_恵u�ŗh�M>���&	���
�Ma�3a@EJ4U�	pn�QiBd@�Fnf������)��oq/�X�:��t����S���1�����o�� 0��>y��'T`�z��h����"�����E�Q{<C+�`֎�OF��C�I/]��:sQy�·o�c�>[������ι9�l��o��  ���X���p �x����X,�.O?�^~��׭ҡ�c@0��g�}s���������ӁƯ1��a�Q��������"��G���;�('�P��pf������b@�o��
��'��¾l��Y�uiA�Cz����}�l ��?�x	p��d��p֟�S�'%��G������W��͌lo��Qg��4wb�*X 4�D�'���R���_�}�����@@���9��}� v@��G���ZtE��� �~���V� ���<��C=u�IL�s&�h�����O����eԉ/ }��Ea�ꄘ�"8,��L��/��m�;�;�T���
4P�Y̹:,:�D��:�0V;�؂�q�����cJ�O4`ͽ����;�*�"
(� �D����o�� �w`���h����?�.��q5˭��ӈ(p�B5RR���&�O82�o �y-'d8�i`��O�:���&*f��U}���n_����e��$�@���k�6�̀�5��B7�۲�}F@��7��+&<��nA�8G��=VYw�y�Sm���f.�&y��O����������MJ�b�3������a��LR�ke!�>�lQ[g�;�/�7���J����~| >�n�(e�z��Q5��¬%��Q�1��s�å�]t�}�o����}I\  ��唺/�pm���������ș���?�����_3A�s�2<�4�<V5λ�/ � D���0�(+NL: ��z���� ����4\	i���V2
�ǜ�|��?���J�H��!��A�x��O�Sy��ϕ�f����5��R	���uNc�k����RþeW
�E����?т������RN�����Bä�.���-�@i��h�ij7�l�:��6�����@S��z���s�/�dN5{�&�M�0��ie�)�f!kV�m8���n������r�>���pL碆�=���%[�J8A�4����0"�BX
9�/$R��L�Dc	�*/mW��_*'���B?{�y��8.?���8����KNK[8�c��I?���eo6�EI� �|��@ͨ�lxr m�g�]�����a�a�s�lH�9�#HL�<;~�_Z\�{!�s�� �K�,�I��Ϲ�[��3Ӳ`�Ͱ�Z�e���s����d7�d�������{F�1ɦ��Щ5��Q����̿c��y��:Zp�ߪ��¤ɓ.Zpׂ;��q�)Ù��w�6�ؖL~�R�'fN"~])ˠK8 �q��a��ٿ�]�͇fO,���k�+������Y�0�!��6��5Sq[��@c6*��}b�)o}Ѹ�t�d#͔%k6�I(z	S3(KW.%�xL��^��6Q�VsQ4�ׂ89��3ʩ�.kkH�rBݜ{�xUt �͒�*<D���^[� �  �Y�+%Rm|>���-j���c�Um0��/~�EȬ*%�t�Ȕ��B�t��̱���Z'�jWe����Y攥�.��Z�|��֪]�,�r��k?��1A\$�]���ح��+	�\М������`�_�F�;����4�JUOJ�(_t%�'D�g�M�2MC��؝"o�����^�|�K^iO�F��c�Μfl2�M�}5���˂�Xk3K�a��U[�&�q���������E1w��VN<���6�̉d;3RK(�Y��$U�H�X��E�%�l��Tid������u�����й���F�VQ�8�m��Tm�������Ǝ[�!��	�4zh �V�U��������)>����D?B��¬v/}}�=��A�;���>��7�!�W�����#6'��Bm|��9Pko[���y�@��+,�#1a�+f�k�� R��y�{�5#�a� $<��%�Y��VUJ5K8Lq�ٜ�(e�WT.F��?gn?��iܑ+�dS����շ�dRZ���C��8P�O���@��8��^xi�����Z�ro���ݚj��y��dr�jf6��a�Y�C9f8�����gt�J!㣥4!~�	0*�����͇%F�|`!+��uP��Ϡ�@��_*�a����p){[D�k���ԓ�V�֦t\ȅ�moڠ�|0a�٬C^�	E�0%b�V�l��O��F#ڇ2$��n����%�O�ܼ)A?����2����]ˌ�,��?^3�V�����h-۷v/%N?k��9�� ��w�]��{�}���N����K{{��{��e��Œͺ^��TֱA�J��

�]4��;�R�:������ɫH���l*źb�Tr�a�hݝ���S+���,6߲	y�񚄴%;d�UkBR[\��mE��/Eܨ���c�ir�J�/	_ֻ��6����K�υ\�����.W�'�L����3Q*#񀟌�Dr���t�R���|1T��C��Sh�oξ��B=K!���&\��;�Nf��R2�ZD� �q ��0����Yw�%��Y�J��+b/+����/9��O��yC��_�B�q�R\�똓�|ù?C��ZG��w(g���N��\�=�9��bn8�	H�S�_���޴��#��|*<���}�q:��	���K�6.�tZ�@&��g��U~�Qio�T�ɯ5������No�^{[�>9�F�Y,JM<!��V�={7�䒋�e`&�a����SO��5�����{�m#���J6_�g�yFc�-ӏ�/��6������A���~�3uH��+����d��@Y$�Ql�u;�SW�P<�j��#����	Eb��B�I��IM� ��aɤ�$^�L!+�X��c����A��6*�AK���� ��j�J �2g\Oڅ�U�AM�f\Tyd=�X�o%��B��k�s��À������Q�?k���,4r�܉'*��7fv/�`ʧ��	&��#)���.�0�����=k�Z3������_��SOy�~�!:T�m�j��e�/��!3f�R*ߘ*�_������haT�LGt�W5��9�Ǝ-��8]<h_�(U(d���<%�$�6l��-�ƍ3Zv���t�2e�n2f�x}0����I����9I�[����EL5)����~�#��6-�8Zs�j%V9x[V�t���|ø�J#�;^K �0��X��ĊiɈ�:����W��nA*v�[e��骍Ȕ�M���[`�tە�_^x�����'K�~�9Wˆ� �-��X�o�X�<C�A�`=0椯z6}]���A�@�ˢָo�Ws.�{�t���1״y��1׼�s-���<�߫��P�����|ǯ����|��=��x�;$��X,$˖.�GDk9%;�5󺶾Nv�<UN>�4�y�LIC�f���C��o������=�h�3w��$�mWW��!T��#�K.�PR�.)�R�ʫ�ŋ$�s�(�X�����1ǟ$3f�f	���A`a�7Z�O<���{D&P��/��7߬ܧ��i�Cs�����W��j�_߸^&�oP��D���D$+�LR��V��rӍ�	e�x��g�#;7�(�Z�,%����JqMV3�W�O�GKw|�d£�yY�k哟��$�W�����b� �8���"�|筽g4���Eq>�j�6&����9�~���ܿE�Yč�*�;��<{��A�ܱPp�c�0�F��Aik*���D%���+�ʋ/>/�������b�����%��%'�����Y�����mwܮרV�b���<`R��!�/�lJ^[�P�lX�$�74�:^�Ԥ!ʆ��;���TH����j�Z��#�<��$��D�G ` ��Oa��ú�DYT���+,΋���b,Յ�^{P��x^_șF��& #�M�0n�\����œ�	�%&]͵J��"�L�����K.OrRX�4ΓS���h�q��_��Co��~U A��B��;�����l^���~�����߮�0+��
~���`�E�Yh�i�vߦ)݈������ޤ������n�F	0�ǀ�w�o�Է��<��E�*{�֬�t���.��Ȕ����L�SR��e�ڕ�a�:Y�����N('�C[7wʆ��RW;V�zϹ2k������������s���P���&7\<"���̝��d��#�45�����U2��F$��_��^����%��U�WH6�rE�����eg���D��w��o;^{��`q4A� �l(6)�>�Na$:B뀈"��"��h�9�q0��Zp�ݶp9����1OY������Z�F5���)��/I�8zIB����N�����&���ߓ\�[�Ѹ�i<K�M�-�|t�௢�^yu��[��u�����L�Fƕ
�1? ߂{�|p�U-�
��=���QHe����{)�}�yM�X����	���P��Ox��vO&�8�w W��r�a@���57Ա�I��snj#A�|�+_ѐU�a��?�����ʻ�<��?�S���'7���>&���$Y�f���V�p.$�tNV,o�H�N6nL�1ǝ('��?���^��%��O�o���Gn'�*�O�B6'{�>[���5��꒮���}�rһ��b�G�4��Q@���I��KV�l�t."�W�ʁ�5�y��8���Э�;���A3@ۇ�4��6���
Vv�8},�e.���ð�B B���{���-�&�T�B�����w�!����$!�?��$V�h�E��n���}�����eΜy�ӌ�%O��W���ުm~7���.+�ՐK! ��=4C���R�4������]E�WP���]�#6e9	�4���O�X�A�'�0���<M�)ꏡ\[5�2aPm��ތ�7�f�0�i���s�Y��y���/jH)�$���sP�xAa��p�z�ed�����
��M��Ϗ�J��wW�0a�,]�DR=���LQ^Z�D��'JSS�4L�.W_�q�������X����-�����G,��vz�w�ے���+�
��n��U�R��>������C%����HGgR%,}f[6%��i��N��h��<T�z J����}�Ta�nB8By�L`u6��f�F��z�D�+Ui�V�Tw�F�u�Y��EW����� ��8d��xp��J��qh?G����-�~�
�jK�b!,�PN��E� �o�����wϝ'Sg�&Y/%~p���f�'�lU�i����[=k����W�������@ɞ�Qp��E +��h�*�O^�L�[��� ߄C�1V^v�rJ���E�ʩ���R�-�g��k�Q9����?�i�+ <�[Ț����<Z_�җ4ʏ}�g�}�҈�y���SO> ��L�0V�-_,�T���;�e��ՒN�ds[��������F�+������?����YC#��46~;ٞ�XE��Y3f�G���$�QiٸV�ӯ����p8%�ׯ��֍J1Dc5���)�[$����u�2}�n��O~R��L�u�]��ll&�Y͛7O31�������$n�\�b2��-�8�*��9v���{�:�D�X�����X% ���u���)�>+�ʲ(Gq�Z?�A1.���
�;Ϳ��N������Zy��g�ԝgI��;C��5���6�}���F�G��>������9 �hno����`�?XW<����)|+�5j����JM4Z���T�P��}��0�V( v���j�;������w�Y��'��	�TA�Pv��i4�F�S���6�oʔ)�-W�Z"���>��ݥa�hy}�2I�;u.�+J1&���H�^��9�������_�DM��(��?�ח/���✹s��L��/�W���ҢL���|���H<�h8/�T>ho)�es[����ꦉ��=���5�d��Y��SNx�)2w�\��l����'[l$�8�I���eQ���� �-����Dk��PIh$�;��R!�l�тF�M�O}J��7�������DC���v���$�����rىb���-7h=�p�^N��?���:�������k���Y���n!����X5�j�3�ʱh�PD���|�V5�&��	�ٳg��F4~˲-�N�Ž�ڻ��HM�����)(6vߧ�y�{&��V���*�p� >N_,gzPn��n�����3��g?��ww��SO�Fv�e�����U����Q'.AX�.	�H��69���e�Y�HM]��Q�z�J���y2�gräK�ϟ[���__ح����E]S'����-��!5�<���2vLTZ77K&ө��<�I��d�Ƥ�i�,m���+�Y4���n����o����6.)�d�ZV�ղ)����%nX�E�P�j�x��<����(��s^Uƅ	K�x�.��LP��f��a)�sr�)'No���OL�@$=��&�)��o�;o�A����i�g���H�8�Ԟr��^j����4���L��1�޴ȵ�u���/�Ɂ8�yA#P�� �4?+�փ k�5J^
�4� �|fl����~&�����m�������Z�q�o̲���e��ђ�X4��_���g��ǔ��N��%��l�[6�4���O�|(!�6u���kecK����d��p$"x�O�8��t4A�����_����k�q�G�|@ҩN	�Ҳb�bY۴LB����0ц��	��²is�L�eO9������Z�������i�?� ���E��ԤZ6<����M��$y�:O�R_W���7F��DB�r���fiK[�R�Ԍ��lA�����P$�)鍧�K��;S�uǥ�3R���-���;�'�ߩ3f�_2�i��6C�M��<���8uU�7���c�'���"�L���:媫�ڂK�@8�s�_t�E�\�SM3C�T�4p��N@���~�ܔTF�	�ZQ�G��xs����(<p?|�����%|Yة��T�d��l�{����\z?� 7���ɼZ$�|�C���l��j> ��;���
�Y��"�Բ^
���ջ�n�V
��,[�$;M�.�x�I"r�P�k�dR����'Mn�l�]~2�4�j_�,��y���������)�\V�z���<)���	B"�e�<i���]�!���S�5�
����o~�	o���_ %z��g��X���e�Z�5�bc���J��U�I	'�?�X����
�!g*����"!���:[�q%a��J�q�����~����K/���~�kFr����3.��?�W-�j�<��s���*9LK*����os(k�ݾz����o��,[[*��GT��M�lx�>?4dӢx>P`���_�܁�P�cn�u�*`�Z������`%� 0��iԈj>`e̕�c@��8��s�OV =�q^�!�,ɑ��mfB��"֞�� 2V+��t�2hå}l̾���p/���P����?�Q8�n?߳,`��L��1}����Xs+�.�t�GǬ�%^#uu�d�]��#ߪt���O���n��]�j�W���{�����2|��O�E�`�Q�	چ����>��j�(6���n�g8>���+��( �w���i�(����v�M���ok� �C�fX3�j�OooY�h{i��U1/�HDk�G�Š-ڹ�x)��AP����+�B�h��$H�
V��z��,ި�%���K�mG�Ux@��Mڹ�y��k��Dr�r�-�ӌ騂��2}癚<d���9T����0�PL��'>��>	hWW	.��-
�����@��>p�* �mp��    IDATk��&���7��u��h��#���/V��^Z�p����~��G�g����̾"J��s<[ȭ�B�%�k���?�#t�$S.^�Z)+8̧�|�߄)
������gF�|?sl�c|�#�Ep��1��fT	&��a��B�{3G=Y��~�3�j�ܴ����~�z�Eۣ��+��$��3�h����c,^k�d�Z��駟��k��4���� ���4 "X�x��u��jR��BAM�bT˰����G��Z$�m��R@A-�E������\Ahd?�O���_*Gu�V��������z���yN��M��p�$�����&��j/_�g-SX�4,M�"������ |��!��ZrbEdQo��Z�L������7ARm��ל��@?�1��/|A��=L('����� <��K��I�:Q#,��s��!b���D����b>+��wh�}�@����\rnY�����!���uڃD�g�P���<�W���=�����X�p�V���������ϗL^�\��ˊ�tP��zݖk��|Nj�Q-���~�.�K#-�)��`�B8T�����2��U�����S��4���4�7;�w�v��ш�� ��'N{SK�
�lp� �� �X��}H�k�������v��m|f��� �;��wܡֵ�a�<����r�[,,�
͟(����O5�`��Y����f��v��V<�=> � ZWR�Ǭ�� ��������:JKD�]�|�w��P�
�C��a���Ϳ�#���1�����2��Ĳ�X��e�Y�"�3�m��u�^ܯ�c��]q��p���,�j�8�~40�3�@,�El�j������6ܾ�����I����4&?Wt�xE��=�?�գ��}�A���ϣb�?��(�(�or����F�F�� ��@��}~�NZ4UA��������?c6�Ф��*Y�80�o�k�kXn��?B��g�ؗP��?`Z�6��傈�s�'؀�H����&�/��BIq�Z|�%`]�u�����1c�j���B�h>~���a�U:ۻ��������t�Ι;����k'��Y�.6̀��$eaqF�w��O:7���/	���-|�-��P�;X��@�-���>�C�@؄
p�QI�H�����.4w^�܄�����4�j௙����>�8G�>�������i4Ž��{�/�9|����g�h������_\��v��m|�4���t�w*M⃿s�;%��
6͟=�%C�ǣ�C���?�����/ �|&��M���m("�Ц��1v�V� ʤzJIZji�M���ʭ����b)�7�2*��N^#4ο��d{�r���s�ol��i&��AZ9�ɷ0N��i<��o��,�dq�!��ބ["�z���y���8���P�װ[l��4���?�q�h���p�M���������5ZY�h����\+� J�2��?������Qee�.��(h�O�~}Я�����?��1m�/���"�������1`6��2>ބ�Y�������-�������7�Z^6V�5�r�+ױ����ƹ�?jK&/��&�m���<��o��k����w{�v<��Y��%qY�-t~�>�[A��Q��ĩ�B�9�q�.^���M�/Pp_U���}x�,h��q����ڧ+:]��1�o���i�����RS|MD���$�ֈk�u���LR"���3Գ��7�Ǣ}��њɏA��e��r��ڱQ2P��	U���t�6����iS�6�xߺ�Y�$���ri�����m���9�y�ʼ���{�
V�k��_a�̝ss2�~i%�f�BA�0p�T�຦hT���^��_mCb�
̴R]_/y"��!J��x��L��X\2��d�"�0�D�.@�8�[A������ΔS�}���E�@���h��>��{6.n��z��WK(H�y#���'Ml����`��U+��'#�N��f���LHl���3��k��i5�xȤ����󀳼����m�vaw�]��A��A��A4R���&Acbc��I�Q�`��&%	b����ԥ���l�;;����{��s睻s�.;�J��������k�-�9�9Ϳ����!%�kF}�9>�|QHϿj޼�_�I�%����Fm��%�5á�N�ܔ�ɿ}S�?��6fa)Z@בE�@�,I(Q��H��Gs:�cZO�h�,喖���%ʫP*Z�R5�������Th6]��+������V�v�ε���\�/9|�}F@�n���M�(�v��~}Y�M4�a��Z��V��h� �Ƭ�F��|�
���袋<�h;!��C��j+�o&|xV�}h���F�����^� ��x�o4WR:]	{�4ք�s���;�����O@��Xf7��ȹ���6u�5����%�R�m&uX�Z�l.8�� ��p���eZ[lm�z��h�j��?_1�?�2�P�bs:ϱ����8|Pr��ܣ}����O�������<շ��� �������LE7L�?�>ǏF���u���B��{z�����%�ܾLʎ7��	%��Q\X����FC���9��������8�I��;z�	�����J>�s�x��~��i#��8�CŞ���yS�X���T�/4�UOq�\R��l%��$y�����Z�>K�zp	���A��������ߠue|�AAP��R�j�~S'�%��t�3\�
ȎMm�;֚���v `b��5Η�#�#��N4��*�������3.J��b�wliku�u��Ͽ���xĴ�"���hA�s9�3Np���|���M����#m&6�M@<�����,�ac�h�x�����-����I�!L5�#��*��[X5���+Y�J�}�m�����3�i�Bۉ3�8��r�EV��]�_p���C=�?�Xdn���_�MH�(�E��P�f/�'M>�jDT�X׏�n�{������Xo�C����
��cy�0�^�Sۭ�lh���'2��9��4��E���/�����V�o0��t��5{����ҠK�ġV��q���P~G��b�+�k<�(MχD9Gswm-�,^"�Z��ʹ�{6��įJ!�����]��L.���J�5��H�/UҞLv�)'�e�����3�-�"�'����"�������6���o�Ǎ�}���B�KȺ���M]��KqX*����v��I�Xv�B�u�l:���0�XWZ�)�c/�J���8��ⱎq=�SO�	W�Y6h����x���� "���O�6X�B�|5m���D9(�wSP3��뵃^�*;������L	��=ے��׮��]���߽���x�0k�h�T�|�	�ٕW\��>p�.<��q|yv#Գ��R��/�'��M/���2��V|~�p�1�"�?�"cZAʋK�/�����h�$�G�c�����5ݍ�JH`�C2}ϦS��M}�?�y����4��1���=��Ϝ5���o�����O���Ku��\RB�0;@����o�Cʈ���`1�/n4|
�Qȉ�Ʉ�@M@f<�F�?ׄ�)��v��ϲ9�����Vs�fq�fF���Yw�z�����z��{�����Y{�X�O�y��!;��W�UW_bϳِ!\-ZKe����J��s���iU���W�3�c���t.�B�� @A󧄂�q�#s�5������(�&;X��W_I֬(�p�\@�84�,��]2ӳ#l�7�c#�����*����>��@��G-�O�'l�$�������R0�s-�P	<�/`
�#h�0�ͪzVK3g�x���fq��c[[��f"r�
���a�v�y��C\���t�Ig�t3�����͛�l��LUi4 ��>�!|�{��@�j(e]��ߴ������F��JR<�1{�l���7y�>ז���j���3\qՕV*��b�h��p��d�z����r�Q���5=`�r��U�[� �f���v�yo+��V�T����A��0���Wӓm�u��KLOp�ui���5�`�j ��8�\o������̈�\2�4V��I<�l�/�3~��j��b ����<C��#A*��`�
��8��C<�u��h�D�� �)W��#���O<a+W-�r�j-�4�
ax)��G�q�-�jub����}���/*;Sj����zՁ6iR{�$
�ļ�y��/U���@���뮻|�dV�V5o�6<1�h&D� �|��ޡ�?	;���aƳ�Y���Ѵ��n�lB���>��������L��'���כZ ��
Dۭ\��L��J]I3�U�͛>����L�ٝ�ێ����?�a��L���nV�NVP�����~�%�U�g���0vZ߱,v�}�9}6ָ`�r�r���Z����EK�BG&�;{��9^�eŚ��R�8��c^k��q��M�p�Jh���6))8���k�y������B�`��ϴf�ђ,�$`+�'+fvg���=�kE�Դ�JH��q���/����5�b�`}��}r����͜i�����=�2hȿ��/] h�0�u@���c�Q����3�\��뼪'�%,b����Q����k"ph�'�P59�c-��P��Ѿ!�����nSuJ�ͪ�3+�Ղ��^Ye�b�}�Ϲ� M_�ﶓ+#�[�ol	lP�2#�9�����VjٶֿVB�
�$����,�3A."-?��a/J�b��aQd��5>�	篨(�Y�V6�����7	%�1�|	�gǲ+�{Q���9ԭ 1��׼�Zr���������f*c����,C:CK؜�E��O��Z�iߘ����Z�К�9�v~��;}#��}@�6�LV����㏵r�`��m����k��8y�n!���v�񯱝v��
�Р�ʄt��s]��G��u�8���?{�w1��5���as���FĢa'�X8��gu���6�O��]v�e��?Z�g�j�b�r�\��]�Q^e����͟�J���?{ι��n������V��ץIR�: ����.Vi��c.m�1�����V�t!.�\�k]+XB R�&i��˾�}�q(n������jo� ;�}O�q�o\L�Y4�>�o|�y�˦-C~M~�=�Я�_�<�T��ε�Ge��q��N/R���ݾs˷���V�X�q����z��74�R1^��:�����k��bi�2���X��~�z���V����S��p¤�מj��� ������pg0��'�OO,�R�Y 4p�q�<���G�g��g<�����(�+L	�s��$��IH��ў��
GWlֶ�ؿ|���:"O�5W�\����W��o�w�� �v;g��t�s�5���9�T{F�y�����
�l\�5���㙻?�s�*�k��M�Ԍ^ �Ϛ�?���8� @q,���ԱT����:�q��g����}�����}�q�{��l�vKW
�j�2{�
�5����!�r��'Y��SՌ���cg���aͲe��%	���	�1s�w�z�����O>ڧ�����ο��gҡ�+���;���-�.��yOY_��\�Ժ׮��g@�kw�Zg��e,d�]7��;�Y���ַ�A���B�w��S,, �9?��3������cNqS.�)KRB��#�,q�Ҷ8g��CSH�,�m�N����-�	!��R�Z�U�V{-W\g����߸���m�s:q������sd�R2�[Ç�s�HX͍��
�l���_A_������l ���j���O���O�aq7����D8Wt���P����3��~�;q�����?ֱ�p��ҬH��"�d*W���Ъ�O�V�(����~�"5g�;�Ӭ4�o�}kl�����m��.�e�����T���ݽ�v]���~v������6�c�}�;߱_����'�
�fw��9�����!��������v���K=�e*vם��1Gf}�����g\��j�[�.o,���ڲU�v��'�\��ˤ# ���ڦ�zϸ�hw�Ue�}��x�����{*�&֬�����X>��a�Z�)�-�O��uLF[Iy��ʖ�>˖�Y[e�Yq�}���Y���X���l����
�i���Ӹ�뱗�~�ӱ��Ib�{�i~R�:d>�V�}zZ��W>~2>���W��ǳ�F��Haoq��gu���-$���4z
�3�{�����k�j����7�[�����i`�_|ћ��4�a���3�K�=kJ%,xƏ�㾮��2��㿴�P�͜��=;�i[���{�
u��E�ʴ٪�n;�����ϲt��~��Cv�w��@o���hkuBk��tv�SOO�Ɔ�5��*��]��k�=����k��w�f�q���Ru�E�\_\���A[�d��*��pq����������Gc����8X,��;��}�+�WZ8���ŋ�O�bO��9�6u��<E+(tT��4�X+��Q�f �3,��ђ���Gl��휳��JѲ�!K�z����T�Ǿv���S� ��Yi��W�~ɴO<P�ų�ʈiJM������g��d�>���[���O�����'��-�y�3oФ
z�#��z�OIg8t-��3Xԛ#�^�Bk��b��
�_vɥ����}v����4�~��&��k�-�6Qqt\�b�=���۾��bS�L�矟�ډS�ٜ��y�b-ֽv�v�y��򫭭}�[7}�f[�d�V�o�@fϙ���|��������o�\{��Re[�����e��z��}�յ��z{���U����]��?X�EK��+�;������c�|����BF+�ē�'��{�mT6��O⋇��vl4��Q��{���U��P>�=e�4����Wmr[���!K��<�kš>+�)��\K��������v�G$6BbD�n ��,0��|b�Xf�+�v���RSt��h�/��'��3k��o}�7>G�˗��%�?~�����X�ƲҮ��Z;��|�1o����󛥜�����I��}��uk�zT�BTIY�?��}��i�@��g���{�q{��w��G�	��>���Z���Y�X��O����|�������g���]0|��_��_������HMh���9��?��������Nv�uW��t������)'g�L��?����>�����l��%V�v{qI���+݁��ô}���_Kؒ�/���ooG}��s�9�Ezǝ�s�@5��&����n���8&�%�9kC��p�'�(sV��j��բѰڥJx[&kE���]3�y�b��h����I9d#Rd8HkDZ�f7}9O���F&I:��Yk�e�6z4��6�XJ��v�o�.�x�Y�H��͟��3�я~�Aozӛ�W�j�*��>�яz����>����m��=��o큟�eG~�M���-\�B�0��
Q:�b�>���E��)�G>�	�2y�����׾�5���s#譭����sf$����F�O 6k�v����`�-4#)��}ێz��V�5kWY��5.$hX�b�J�^���dE�q䱮ɠ�,\��#~Xtj�ƽ�T� |��g?���{｡v~�����?��c��@�r�nC���%� �8�˰��L��28d9��V��{���� ��A���}�a���w �7��J���d}lrix<�k`ԉ���l#P�(X�P5dU�Ҋ�c�?~z���������� �F�O�s�y��Y�{���_��g��P�(r�]v�;�|?�����O�����U���w��{�lmm-�l����'!�<b�Z���t��s�}�ʫ��z����^�%'�JK��Ϛ1���n��k���'��L�omi���n����暫l�=w7��#�����Qجh]���W�T,�C<��s�z]��YW���~�����;�?��O4��tLS�s��n���������8�R�c�m�m�Qj����Kg���њ��gCW,GR�ӡcX1]���,%�	�䟁2���ޗ0H�x���@'p�c��lL��
(    IDAT�?�K��(IP58}��f���۴i��+�� �i�8^g��e
�D��p�^~�e��>��5�>�����C=�� �����<��`�|������ͯ���cOe=�z��d�
�Z���/��?�Ֆ˶;�t��_�tv��CMY*�<s֌+o����N@����ϤP��M�o��k��%m��?c^��&Y�R�����1�%˺l�=��#�<�@L0Q"�/���F �����O��a2zz�{�v���/Lڗ��I�Q^>!d�V�+��P�V
OQ�7�T&e�T�J��-�.g=s��?)�7raK�'{m�[�v/�:�B]% ������Fxr��(�F��;��ֈ�C�� �G�����-���W�"<�M������W�}~G��-Ͼ�� ����:�i����V�E�����˭l%k�d������)7c��csm�=��O>Ͳ�V��l��η=wH�ӈ�JJ:_uǭ�~e��ء�$y)
I~������ra�Vu-��}�y���?�×�a3��̘1�Nx͉����y�;��mh�Lc���=���k5u�5�M����s��Ga�,.%em�8�-��]8UCMO���:�4 w�d���0%����2�!]	UC�-���U��� Ц`3�x%��Y�>�^����7�w���h�?�n�Z9
�e������{�5׸U���8�������> w�ֶӦ{�t
5����ş�/��gS�~A��;ﴃeR%[��E����l� �@w���[�~�Pr%e���n��ez�m��Lo+:w�\��׿�B�YT�����O�{��n��KG��BU�C>8Ak�Y{G�
�6�3������h��Z<�v�a'g�;&Mqg��������}4�~����JO� m�����;(����3�BMSZ�c�+N�x�>���f�j�rմe�L�R�lE��+�%}z��L�J�@-\tʇۖ�!Z��X����q|�?�S��ڐ��8|�͛WK��8�4���]w��0_(\�3ڇ{�\[;����+.�k�X���G�M��߃F����[
����>$�N�h�\.c˖,�����}�����w�o�Wڱ�g��S���6~�B͠�R3Z�B�����n��扨�&��~g#�'��5�J��\��:�.��"kk%��6���`)0�CC�E��~�Y������MQ�C3!i���������'�͉G�$i�\��@ �s����e�� ;��sN��g��-!]8`d��cx<�f�kc��|��˄0OYX�ކ-��Sx<�����7Y+q�'mN�$И�Q��Q��X��v��w�Ã)ثh�(a8|k�S�u�a�0c�������l�#��Ѓ���q��5�чɞ'a��5�F��cO>�d;�3\9t�X.c==y���m7é�.ϱ��ߙ|#��p�w�(����5���sN����w4mve��7���W��N?�4�o�}|�x�\��0���g?�(����9*�8d�}�;���w�B�D� B��n�{đ�+��	5�N��6!B"u���8�{�>��zp��h�bn��]�A�(�{0�C�q�x���E��C5��y��������|�=
�9߬m�c�B4U(�~��b�ࠏ?�S�[�M���:1YS�t�]p��3N����˗���w�=����/ae��^�����l~�����ӿ̐�s@d@�f�{5ΤP$Q=$xQ�
�5a�� PQ�
�i���%��jqL��S�AN�Ϣ��f���f%��d&�Ae��H	#������R3��I�fB��_��q���7�x�GQ'\?���ˎ;�8��ǧ>�)�&eQ(���I���j�����{͝�WX7�^������K��i��B6��c�?�9��W�P"XZ&?E�H�H�h�7��?�X|�T��k�w�fD��b%�ȐEA��T%�ap���KfS'O���V(B���ڵ���z8w|�����w�?�������0gP:�~�pSwE��3X��@�?ɠ;�s�?ȸ`Q<�����\����, dBs��s:�Н�_Ӑ�I��2�Z�L�6�IP�1���D�9L��E��R������{,�!�����D;xꩧ�+$���U�g3��lsn�|ˎ�4j6�ֈX'�
bwGwRwF�z�IO-�=��r��H�DY:^חe����P�?�u��x�Մ/��!*����N���1|�����M|(� �Bӥ\k�gl�L/��a��R���P��U6�����w� ���W���܅	<K=hk�@�ȳ�?��FB: c�τ��sf���K�O����1���dVk3q\\S�8h8C�I��\ t&�s9����`
@����4:i�ٜ[�ݲ#�<K��Se�e����ޱ&)������� i��ט=�u�{�4O�?���xF���El��'�7 �Eϥ����R);�f�I
�Rb�^�ʞ� 䂕��A\K�B��<#�f��c��N^P?�>��k�P8��b:NV"��t����*�^o�qo	�۪���zgwv�G�'U#�_�Y�˱V���:���L���f�5_���ٛ��f�����X0�zg�y�Kw"pTq�"�bw<�s�[vb͌y��-��ZІw帎��i�zz��@����k��aL�H`p=S���@?J�ñ��艐 H<�8�`�q�(:=��%z�����e�och���I��TEb�h���/A���~'YiB̕�Z��,v�B�� ᭆJ� ����@�q�-��c�T����9�������|��F��+��A����8�J����-���\p����U��9oٲeN� �!�.Ƶ)���q�18�ڪ��,�X��Ġ\oQp��W�Xv-7)A�/kU��h��2؎k����^8S�����?9��e�d, ���N2Syf(�M3�SVl���%tmů����E#�ߟY���3�z�į"!.a,� ?��\����%@�@�1�<�����K44�+bc��j�R�5c�U4�s�����+�����$ˤ�yZ��Fc��i9G|?�7�o 2��<��^d�����Ƶ����t�s���L��?~js�4O=
�+������
����c7��c�����$\{C͸�Wq@��_�[5�O@[��="K�-�t.�P
NU*߃�	n���H�}�e�fp'�[a(���A�j�["��'��MLw���O�_�g�/xA��V�ϱ~�Jh�M�=�;��'�{�ܱf�9k�շ�r�M������9��Λ{��7�Xï�~bs-6W� P���4����z�������2�!��Ŝ�Kۖ[��C��@JA#��M�	L�f���a�|�$J� 䑲�7�.��2�Kg(^�=���@��R&��c�C��P*�|3k�3�y."Ɉ�"�&�l�X)�G�Z����˂�r�eE�;�b���.1:�g2D�T��	�-������U�����������a�$�Q&�%uJ��p�4w)�RP
�R*bZQX bc�Z�VgΚqՄ��sf%�﹬����I�b�I+��%�%�X�/�q}���LҖ:FZ�6�ứ��� ��5�`��e�b�S$[j�{]�Q��1H�;�����k�}��k�����o�|�����p�KQ2^ԣ�40׺�K줓Nr ���?�$3�9AԒ�o��,$� ��K/�ԭ	���.S$���p}�x�l��WG_�E��T YB�d.��2XE��Z=z�(DT�0#�.Z����fB^����ɐ�V�G�Y��=�St�ش�x׎Ώ�0�;j%D86���SF7	�f�w+������6��ɒi%@�F�F҄���8@ I��uo��ב	-gd�o��&�Hi2����^��I0ΓbPԥb�/��͌��o��o\;�j+N~4�v��������!�4.�2 ���_���[n���Ϗ���	'��?�>��>H� u���E� ���p�O�k�B%YƙZ7�?k�+�&�LLKĜ����α�pl�O{q?��P�)����$�>]�L���P��l]W�RI�j���V"O �V[���L����������>�q.�D�
ԳC� ��19��=�QH���o�1標���My�c�&K��)��n�$��H���Ц_AIk,8q�rR�f)��j�~��Ό�ų�ŕ�"��b�������B���ȣ���[G�Gk�}>'A�"f�iA�@Fc���/�Ў?�x��hŃ@��T傡���}��j�r@�0�\�gĪ �\�k�h掁�@�� �i��Z�B�2�����
1�N}��A��k�b�\R�����O�aKD*�%$ejs9B�O[K��9�J�leچf�ҫ�}(�b8�w��>7e=�t����E!庶�:�M��Jоe�H�7��'��ߌ�g�\�M)�C1�|�{r�2��M6�&De���MY4�����G3�5Y:��M��^Z���2XEn�`���_�4�XS��>����$���_�����������?� ^P6��������~F��: ��H�BB|�_p����x�8�K"!��x!<�}xA3Q�W~$i�γG�/��WrO��O �Bk�H 8��K�-Yh��͍Rj43��y����'0K!n�+�)�y��J�`�,��RVJ����)���Vk�%m���-�
���rnsC�s���hj�Y�(D��f�'�\&`a��Λ�=��7���1��] /
��/N��z �OR\[�!phf�5���~΂���#-8������^,t M\&�g�ӟ�4l����e�������C�w�ԃ�'�ZOh�O>������
��K�U���hd�}������՟�ٟ�` �n?�n�kB��~���=a�5�r��w������G<;U.���K�q�G��1���=��8���m��b���L�c!�fU�y��UI�80���2N	��%�[�q��L%k-�i+W
V�!KUKVv�?g�
I ��M��$�������]{�uȍDM)@@J�h�P�"D
���w�ڷ͒�"���?g�PO9[Ўpx[�qlB"7(� x��is0DV��c#��2ɘ�\�SE��h��=�G�}��~#���黥5YL�hƸP헱!����g,�k�Y���a��)����:��g� ܧ�z��J�_�0������q,V�b_�tVׄʁRB�#נ�V�@2�9�nR�@<� E�i��\-���W���شO=�C�S>p�Y|���U�k�Vm��w�=����V�B�bm�f��Y;%*I�*K�:�g��a�w(/���=g]��XO����2��;d�y�1+.�D  8?q��2va��M�3�q�C���O�	�GYh���~�8�B���0���L��Ϙ9�	�̥Y��(&II4H_6ٹ�ז� Px�����pP��<��.���¡x�E�L#8�-�x˄	�F���_^�/�;�28cΟ���
\��g�6�r�\1��5'�Ua3�����%*ǠBݯT� ��b�E5ȹ����|�r*� �i���7���Z�f�U���Z��O;��8�Dˤ����Ҷ�������3@\�;��mP'h�:q�А�,S����u����ڊ]�կ�j]+��Zmw�'§�D�T�X����Ж����c�r	氖���'�x�+�̹B`����Q؍a(��1}�hMh�oV�G`��
��s�:�N8�P��2���n�ZK���|�,��utLu��{���2��Ln3�̖>���駟��R, w��WOc�_�U�P��Sc/�L �����e,�{�t��
�Sē@_}�.�Q\��=�� 8K��zNC&�8BD��d�i�şK�������_�Z�c[��5�nf2U˦�V.��i'c�{�IV*�[*M�i�Ǟ���@��5�O��Rٜ�R-6T*�50�+�T�h�){��Y��+�h����k��?��m�]��J�^�)�9��4�VHyd�Lr<�p�y	N�W��?����;��k�S�T�U�,m�&4�7��$��*!��s;��o��P�![�b�����قE�\.��D�;��C�SN���lk�v�B��tcΎM$�_�_ٿ΅��A��sbPP�q3���P>g�vz��{�s���|�Z�W��}B��?�K
@����]*�������6�4j�6'?���:�F/͚��lTzAsͺ��(�4u�g���/����@kF��^ti���(�_�g$� A"Kgx�|=#�'h��n �{���٩'m�j?�>���l�v���<CJ�t��Z�m��1�Z�H-�ݷ��Y�n��"�m��Gm�o��RC�*g���h���w,ߛ���Z��=���J���-Mt���[�i�C��d���Bi��j�+�B����ʷ_a���a��y��.��ϡ�at����;V`�����#�w�Cה�P��'4�7��_�(��g߽�?��&Mn��U�����Gg��5�kQ1LJ�[�v��Î��:�'��&�0>%6q<�t��ALv'-��@m&mQ��EM!d����أ'�V:p�4,�x����	��T��c	2�
���" �!�/@�˺�8]WB�ϤM*�?��ba�k5��e��Z��H8�&�6���&`��1#��!�3�ϡ�U���~�s�k�ԓ^m�r�����mmڶ;��`ي��M���e�mV,T����1c�M������P���gh͵Y��gK�κ�.�j��ҩ�u��ؗo����X�rV&��7��g���X�g<'�G�[Y� �A�-`]��>�(��u�㼟5c;kɘ�p|rr�Z���Ckٌm��L{͉����z�C_p��9Y��Yi�����|���F�>���ʦ�6{��v�i����=��k���^m^x�z{{<b�D��F*e�Ww���C6u���_��ӎ	��~DgP���#D���	Ĺ��o~�I8����I�
����ϕ���S+������|ST�P��w�ѵ��w��a`�������@1S8fY��.Y /�'*�*�����
J�=�/��"
(~6	.�d�����xw���NT��e3��}�k����J��*Ռ��v�Y;�DҥlҤ)�΄օ8|{{��\�����v�P �{lh�ZrE�Z1���4�c)k��]f7}�[��b�T�U2P��T! 4t��=6��Y/�5�
�V^���}���3J�J�s�8�^RV���.[��{�鹶�7�t�?T,��@�֮[o�춧�~���ʹm=��[o�x XF�O'y��}b�z6�͔I���iӷ��2���w�=��+v�R��-z��}\S��ށA�Z�e�r�-�׽�ӳ5�8���-��ވ� �����pCy�������/x���!�|,ir,����j�c���Oc.���{hl>i��$��<v�BH���c*�O�P�S�0�"�!v��z�N��K� �yLO�7�*�/��{Z���;#g�$�3���<�4E�o�R�>{����I�=���>�fZ�c�^��nX[K��������R��P���´��&O�/�io)YO�E��/5+�[&�f+��K7�a��a��"�ԁ��y�u�A	c\Q���%������2��>����m�f�>�kKY�e�[�x�w9�500d�m�mɒ����V�Yo�\v�t�V,V����[n���h���&4�7��K�1lםw������X�w3�?�y����c\SX�|�5Pu�?���/\l}�f�W��~�b�z׻  z���Hh�LL6� �٘�9��u�U�\킀�!�nEn����8uƂ���?6�v��f�c�޹��6�w�99J�Ҧ 8�x��f��`9�b�&���u�����t��9c���Ɗ�QB1m#��A4�^]�T+���X�H�q�;�3�v�%{%Zt-����
���N������'a�r�U���.Gٔmw���oZ��B�J���th(OC����X�0��{��Y����׻�o�d+���7�ak֕\�SF�	�    IDAT�����_�>ߓg`�E0�\�`�PY�ˏ�dt3�(x0X�KϷ_?��}�����Y��s�u�;x��l�=�س��vؚ�}�������v�k�+W��<�ŋzm��"�W���s���lOw��F���Z.�>{�e�|�u�Mm�������c�y�ў��l�"����	�d�֓�%K�Y��j������~�����v !�����y����L����H<�y��>��x�v0�C�9��scC��[��r�4"J�F��{��>��̝�hb*@�W�t2_
	i�Ҩ9^��|��/��:�,��U��}E=��~=��Gk��R%(�N��_^1=U�p+%IЮ��Y �h�T�:�9�N<�(�z�Tm�=�:�Z�gY��/:��	`$w��������� ��YOOޓq�����Ֆ�-�j���{�k߸��v��b��MLmE�RԍVI<���d=u�Q��o��6/����C^y�^}�}��f�n%�Ս"8�����_�mGq�M�:ٞa��*EwDS�(��g/.Xj��$[ݵ�֬�O��=J�ZM���{���|<�-�a%`��o������c{���X.]�%K_�_��#;����R�ŋ�@G�˶8߿h���ڳ/���~�Wgd�����?\�h��ꪫ<��+�q~��pΟ"]J�  �(�J�l���q�V��ǠG4�Nr��$��o�� �l$H�o,�w�e����˚a��S�� ]O���|�)��m��@�?q�|VuZ��)�ɲ��� _����	�RB���[b!��#�w���W!�
��5�,U7�v��N�לp��J�VI����l��if���0�=X�sV����RgK�����2x����P/��
C�V�H\%m˖���[�ۖ-ﮁ����o�F�����b���_�c��O~��W�r8�x���|�#���z �������~�=;�l���J�h�\������-���Yת^�d��>�i++V)��ӟ��-\�|�*���X9���\�p�V1C�Y3���|��V)z&�7�q�w����UK�o}o����D^�p��*-�pi�~�1^G�����(�t��l6x`�Wac����Ss�=6��Hӓ8h۪�7����? ��;@2wp�l�_��מm)�Z!���UV��b����/�ιd��X����,rBD������B8��X��Q X[��v�\��ƽ�YOj��#Z��F����G���R��R�;o�T�,�1�Q��]��l������9�
C��ɶ۔�{Y*=9������\�t�ޝ���{�X9+���0���a�������
�P�ǭ��B��5��ׇ�|Ya����{��w�XSO	
������^W��f�c��"�W�Xh���ǎ�Î3l��'j��Ht˶�ܧ�Y�J��m��N�go�¦M�i]]��N^�腭��h
�L�J��I�f�d��Km��w��\������Ͼ{�`��]���4����x�R��Zo��%{Ӆou�`C0�ԭQ�8����cs:/�¹3��h��).��7��V�o��f�% H7��T�C=T�×FkYr�rGE�����
@0 ZD�!���zj�E`��gb>w�K�)�A�?k�{B'��  ��L���r"J@�kp�]w���p-��~yQ/�u�f+�(4{ u�_JX������W*���%����jf��b���#Z����ed)���@��U���r[�R��[*I����c�D�� 0N15w�Eفh�W嵳P ?����R���B́�&��ŖIlĽk�&������18:�l��նx�*��ڜ�7�QGo�t��>���緿S��}��U=u�J�&��3O�׿�4*���}���l�e���L*k�\���Zg+��m���|��j-����"�ŵN9���j��{�q��a�c�N��x��s����#(-Sa�lZJ{ �R!�����<�N�����bߍ��f��W	��:�ی ��Z9�ro9��q��g���# }��|�߬)�G�>פ�3k�sE��i+�D�EMd\�H��C�C�1]�G�����p�|�G+/�<>�R��M����J���H����B�E%�s ��f�3BI��uPM	�I"��$y�9GFio��G�n���<R�A@q����q�E�\��o�r+��.�[e�kW���-זAY�5k�=}�1y���^o]��-��oo~�%�݌�\J��w|�~����5Дc���������[�\�?�r������9�_����6�×����O�`���ˎv��o��ӦX�2d��=��Þ���i���l۩����w��;ʆ
%��@3d�C�F0��DBew٤�+N��墕�!���G����?����3��(hȊ�Q��;�K\U1���#iD1���hq��@������ơ m�K���h��%A=)	`�U�
�qM�����x�y���`�p" ��{�zR���� �zQ#	3W�+������'Y���ݳ5*��y�н�
hᐸ݆'
�L% �?k�U:C�^A�'1ܴ%� �u��ט�g}0�c,E�$OB�����c0�(x�;��x㍶��)�^�d�-x�9[�b���-ז�l*k�C�6y�6��:�;�H���N��jU��t�Ͷj�jǯ���`fwv~3ߓk�hB7����N���>�.��ki�X�z+�����'6�U�8x�A�ٱ��i礡�~;X�s���J�\B����4O{�����'_G�� [���S�WR�X�������U2��#�H��[���}x`�`�5��.?�/-PU,9� �@q,稜8�����Y[�8��(%\+Dk��*��{��f]J J���)��
urj��֨k�������Oi0�.Y�5���(Y����ܡ����h֠Jl]���U16�����7�D��+�(g�X� ���1���1c�Q
����lp`��Lj�+���w�e�}yW��:m��6u�t;���m�]����^f��q������En�F�?g��������S0C%�8��'���:�u6���z{�[kKp�6X6ko�_�Y_���P��~�;U�A�x*��BaC�,��niܿ�6�2/�H�M [��9�3�w�^�:Ná�V*��ŝ˪�󷦕FmE��7���}� �F�����UF'Bց�����u���@����7@3�:rfs�"~���q>���ǰ�P�$X}���.r�A.��i��qkP��AH{�ɰu�ţ����M\���o�;�� �[7RR�sr���Wj�FM�4X&��J�HI���t	�ׇ~�)�%@��B@��(��ߡ�O?�u64H�G�r-T~�vE��E��nc;ﴫ
���p�i�{��ahO�I[�H�k�WR�ab�>�;;���ɿ��.6}�v�h�y�v�i'������!U�g" 6�SO=�� ~O?O��)ڇ��?�����W�£X@d������
4I( 4:O|�V����<q��`ߏ��=+�s3�6���%�� ��ﰒ�S�$��|B �D�p/�s� 7���zA0�9��>` �1ψf	�@ @'r,4��s��\�Ǳ�[օ ]��m�X�xP2�څʀ�E&?	��9�j�2��ƥ��$�zR8w����	�>��B�}���������哀���� M���>hN!!,K�qf?3�8��8�o�� 3?*���>��{��z<(ԛ��z�ɧ���g;�8��|̳��|���}�1i�Sy��|�������Γpk�ʷ�C�'K18�B�謥� Tڴ�^g������Kd{xm�G����9�=�����#:�J�|1� <�lhLB6�/���������9�n��?�(ʹ*�K�s42�wM�R��ߥS��U`���%��a�3�̭Z�1�k����3� ���h�h�QQ�P�3����7�FP��$�?��5���M&J���V3��Ij��+!�)���q\g��c�<)����M��Ki��s�GO�I9�c9��4�kS�f��u��(��o��M4��$%�k��օ�O~��v�]w�~���+Y�{V����gM�A	P>�"�v�q{;��cm���9�-%�2tt��=��S^.~ͺ���*�vL	��dF7��gΚq���~S�q��s�t~�'��htͿ���R��b�r�!�'�=��͂$n�P�+�8������C(�����a���� �Kj7�=4�K.�������%{lb*�[aS�V�{�D�H&|�xw����"`�?��^�Xjr�h���������@փB|�+*��կU{L;q�k���N"����*�W�e���RX$|�'X<	�'�S��寪Y9��y�������0�k�W��^�`��0��2ou|-��F-�3�{l%�<f��|�U"�'^'�k2uk"~�v��; ��׾֕;4*��ЩJjd vS*>�
��P<4���|~�uw��|�$	��o�R[[(3aqo�Q�����C�XXmI|�����n�9fk�xQq��c�ɇ2@�3���dx>��N]s�5�9�}��j��7׊�!XDlLg@��������29�1�[m��ix��f�% d�|�S�rK�Yw�$?%�c��p��E}��qȋ�q�^��ω鎀�8�Ѓ!�������6�~|l
��>r�J��X��1��V��յ�@��f>��H�c�%��أ�:�kn!9�%P`В#�?���<QK�a��k�BeCoK�w�]F]\�}��KC�N���t������S�=����'���E�/�G�F��<jxѲs�׆j��˨�<��4�S �w欙WOH�������{.l���}#0LƆQ	A�	�b�VE|8Y�4�V$��=I��?�s/��v�2��Фah��Ѧ�
8��B;}���~����}�V�lGi����Р�0Nd�G[4��� x6At��8�3��˓���Q��J�s���$F��s��Xq�����߯��$�����f���b�������D��3vs.kF��a�0��^z|N�L�� �5Ф���y,(�^@>^�̔�4p�Ԭ�@Ŗ����)f��P�m���9�=��W���$5�j͉�1V@��/��-��ZK�
�|L��~�(���u�?�/��{Ml���%ߓSc�	>��l��R5�lD�Ol���i�M�?N36p~,���ȩ��� G�L{q����Eb
a���"�t4&(�[��-�������8xd�5Z�5z	E���B>c#�̜�<p�18�2!��)�'�G��<v��3L~��㇫e>��蚪���̋gB� (P�����<�� ��j��<E����B�9�lt*jJI�y��x&	]Yc���"�D=%eFV!�s�@"`�.���l�40��1|ox��Эk<�Ϲr�K�I�3ỏ,(~���o�A c��FBIyc��U�c|f��	���,�$�����w�ynRKsd���]M��9*-K� O�F��C{h�j�)Z��Y����{�:�+j���F}��^2�"P�[���E��O�<�|U"�K��><�B$�k��]V  �s���K��gNI(㧴a���9����"�T:��	8@�8��?I�=q�a"���z�B�)K��~�[���Nn��-�z%×h~P���Pn4�MDՉ�A`IS��r�+p��\�����O���Xh.CUP�:��Q*&�w5=���i7����+ƞ��	sc����x���6���k��fb�'0�"U��T��C�Ģ�糁y����)h]C�����1l�Z�i"h��67��Xm�,
QͿV#q��Y]�.�q/�+ A�:cD������.���g^T�pt�o6�cO/�7O�J�:J�����	o���d����Љ����Wq�����6�����B��f��y.��uyv :�s�.��_~i�Ϻ�'M�x�y��K�9�Mx�����j���P~g��x.��b�C�I�"��zI�F*ž��y����8]��>ße��Ev�-��s��4��p�&���ԯ����#+T4m}C�F����'�7���Fm��i�	���8�e����E68P�����j�-Pa�0@4%�H��8�
w��y�������/oX�Ζ�����$����d��Ҥ���pH����qrj��\[N]�<7��	ϕ0�W�) �f̵ J��$.Yrr��LkO݋��YJ�R�g	<���@�����}xO<;�������d�] �:Áy�A����ȓ�@�B�q.�o�w�8i�|/�Cd2š�Z�::s�G��"p��-�_*�C���}�(����3O�z\���W�%���4N
`.D5SNF 
5�^�~�
�1���wD��(�A����h�A&���K�!h�ld5��si�V��1��,l4=ř�@���V્΢��rP�D�/�7�m��N�F��ܺ�k��ъ����_��X����c��>�y�<�( �U�8D��&����̭曹��&�Gh�P9
��oU�Dx ᙹ'�����e��s:R*��15%+�u���R3���|b��L3�C��,7�A�<����^�7[�zUT	7D�[ �Q#Ifq�ŦM�nm�>��W��/��^*ݩ<��o��/�#���=}&z/����b!!�b�<c,0�	�f�~Bk�c��7�z]C)[� �5��Y��@�4|i��6��r�rY ǰ��81�R{��K� &��.�f�� ���t�fZ�,�!@	s>�	����|��4n�A�.m�EEc^x�>
I߇����?~�[J����o t�K������;2����X����,XB�S�>�g�����EY(�RJ �
�s�hA�N��O����`=���f���F�'` I�c>�`��#T�>=!�*�)8��Җ��l֬�m�?�Ψ����CJ0�D���t�8�'"�_B_�@���W�ޯ��	��[���sD���#��3g͸rb�z6)�6q��e-�ZN�@ҦT����X�\O{�簨��T�M���a6�;��@1�2'��M!}'͟��YX�i���኱�"EkH��Oir���U$��;]W�%�CTB�T�ȱ�N\�8%����Xm"}���T=�EK��E;4N\Ka|�uUs߿��Dhh��H�_Y�������xZ���3�|�s���y�=.��g ;B*	���yF5o��ǪDH�"+ �
���!�<3>�I���M��g��)�Ce�1��\b��GF,%O��޽��U��Ο}Ʋ�S4��a�n�������-_��È��?/�j*��p��֐�{	I	,�X�|m$ٕC���=*�r<�+�=���`�(	o��Em������v�Z@����`�y�v�I!:�J�k�V[Oo�ggs�����]� ����=Ĝ�&[�D�B� �-.���Х�iaJi��ڸ�X4A��:_Z����o�K�u=	�%=���_�a�kSmI�g\��3��c!!��g��������7��q����8t���ԙw��́"� w���#׵��3]	@�g�p��x�N��ܗ1�;�y\�.^�[�B3�;x>@��Pj���0� @�X��VD���
5��9�Ѓ�"o���5��D	8�6B�p������h���RY���5��/<��e8l�����<)r�'��%�N��qh��E�tl.�q���d<j�Ak��N���'�n,0�5�1K:�O��ϔ)!�pg`��AK;�������B�z�lhpО�;��1[�l�ku
��s&��?J��̣.���"b����\��h���c ��౳Y�4���-�A֎61 %kF1�S��H ļ��@�1�Z	��'�%�_�Z�w(������[C7�p|r�z��H 0l~QE\S@��XY<��=�9�q��:1�$�Psm>WY*�z    IDATG���{�
�^d������r�yzO�{��Eiq�rR���֐��|�;�i�|�V.�?��*[��n|����Y�~�lR�?~��n������~'���e݋��w�:s.g�[#IiW����X�d�c�M�����[���γ��	߇	��������������s;����_"G�4L-D��������4�a8��C��K�l)i�yY��i{q���/~�i��f�$�� 	��l^6*��hhp�t���'�$j��C�F��~i%��ka��9Oe$TZZT�֭�$�44rT�P��Q�]�s��X�m*�I�%�7��g���6�(�ሿ���2�f���ҸD�	����%�%,W�Y�þ��h ��<���`���@�7�Q�9�&s�0S�/�Pv|^�!���Hg:��k�tnSN;��3N���/a��J��(Mc�5nex�V!�Z���:��J�OL���)�-L�@N��E�*a�g�k�0�<� ��|��x�=QVX����9���;����K�ٝ��/W )c�أT��n���s;o�i��15&�EO���k�w���� �k�Hb^hlm�9+P�m���Z�}{��&d�����}�Cd��qt������I���
`�|�1�C(� uxӄ�Ȣ��8Wi��% `�'ϮD��;A�NDY+�4cA��&Y�L�"ekSIK��-�������L*8�Ѩ�bQ�A�4�ҋ���\BUVS���$ 4��?:���I�g�5M	%���<�E�i���!�_V�)O|���xM�9�N�_����GZqpȆ��e	�N}�j��p-�c�whiks�v�i~.�>p� g@��s�~���}$|e��j|�\%<�ȘB����y������,��T�M,L��BHպ��ح��ns�>�nO�k٪�7��:�t~�;�����ς����3N;�.����Q�`C�}�����?u3��6}�ǃ��Cl���I�C&�x	�㚢C(`�$#͗ʞPI4{x��_�E�ЬT$�x�����$-� �+��&���*G����Ǳ,T�?r�/�C�ݠ�dxg /��4�wBy):������f���{�]J���%i��1"��R
�$�%4e��/1� P�ঐI�ב��8�l�(M_օ�Be1�>��/IIF�3��
VF-���-?�,>�S����:V	d�{�Æ�/�u��3���.��?�iT��tu��=�(e��^Ƶ�oPl1奧YcJ�"�������z�2��;���D��ڿ�Jnd�xF��`~(��7_dS&wXGG��9���#�sK���
;�#m��l��P��>���ZWW�_��i2����3���|�Ս��X�l�]w�ٮ��Z�2u���d����<�+[�n��n���f���vԱ�ٌ�;��S���;�9~�T$��� �f�V �y������W�8�BZ��IҒ�*s\tE@�pB5�fA�*U�J2c��3�8�s��� @������Y���L[�c��Q�%pR2�l~� 'c��R�8�oi�G /�� ����ǪSct	'#�~��$��;q�S�=��+��se��)*��ay����D�`n%�@�DH3�Ж�Tm Y�(i��ro��i0���ޑ�QLX�N�̏��1�'��e%�]Y7D����;�_���w���e�"o�@�&��Y��).^�eoi�GQl��0��'ƛ�ZI�i)����m?s^=�Y��~���z����8�;�'�:�̳�^�T���h7��U_͒$'t�������{��6��-�gLJ����O�޽��=��\[�����`��q�-����U�l�̽���Z5	 �� ��(��g_�j�0�p�X �����E"ڠ�O(��Y��}Y4lp@P�,N4o>�"�cC
X ��h+���V	�(-�c�X��!�@)^�s���@ı,r��x>�%@����#��Cyj���A��{S�Ǽ6�(t# L?��H(�
!� 楱`��L���C��Q�r�ATcƘ2�*Ɔ�e�'�n�B���I�$�D�����q��K�zi�+	�f���X!��K�j���lHn+�J~����4��������ʅmʂc~�����Ip��!�G`̭, �7�Ǿ�={�����Z�E_�'�>�}A&Mj�� ���i��������v�gy�����q���zH�VͿ�̞3�������?�&ɤ�ɮ�Ϙ���������]w�e��l��EV(�ͧh�ۇU�cU[�v��=/��4��6��j�ڋ8r�E�_�$���~^r>k���=�� �?]����\� �hҮ�[� ���D�R!�A�@6 �6�|/��84��4{�� dXPb
��9;ƞ"� ^X�S[�����pGp�Mw�N^7��s�cm>�͙c�X ��+~zG�LƵDQ-�=��8�ZB�p��5�ye�r�1��!�$A]��;z�.���X��C�^� -
e��7�x��h��2#5b�t�Kb��\�ԓײ����y]�J�p]E�q���z��}]?��5�=뚦8L���/� ��Ų+�m����@����xɋVA�kZ�RM��E+��l��e���o����ו�{�C�6#�3ʺ�`���ȴ���OHh�]��?�{�*%�f*������t�1V.��E���\�i[���V�\g�b�.[gx�;rj������,�йP�3�I�������<�T�qj����7�KCf1�)�bt R� �~�3A4n�h@y@����;�	���U5ZK+���}i��>���3��{��#\�c�5[���ϳk�а��F�g\����b��������v���:4�l�XQ� �;Vt����M��jn��-?Ϡ"p��^ ��h�oE���s�K��N�g�o�%̽�L��M{�S+o �y_��~1t�
�y�.`d�# ���
�'%��[ ���Qx��|w,����σ:XÊ��3����}���`�ux��3ԟ�_��m�ݶ�i�;�g���"����\���y��*�zM���>��K.u*k��.o�l��Zص&����	M�t���\w>��F�?���g�W�{nx7K�.�g?���䓏�je�V�Zl�{�C͕T��u�ڲ�]68d�t���+��pL�����ᣄ���S� `Cv�a.���tg�Lhmti��4mD	iʘ� ��� 0c� ���f( �}�'��Nc��A��u�h��f)��}�B��0���1B0�q��b�Z�}b�I��-� ���(ʉ����k�D�W@�� ��;B� ߈�r�s)�|��=� c0�Z<'Y���.��� o���%�'�P�=��C���R�����o&b������{���w��?��2����p4�{��c�QV���>�яگ~����e�w� hտ�˿�� ��1��S��<�����;�C��Y�O�y����\���6�_�g�Y`����.��N�����������������hNa�U�o��Wv�y7{�{n�L�b^|�~�����c�R�׺V/����\��n]�-_F��6{a�:;�����x�ob6%�ڕYy�%�x/� �x�|h����O~�V��E�H!~ ���E�p=��j�9*��DE�<p��@y��@Bh�@(��P:�g@sAh���Z�|T����#@u�<��=��=TE��Z���O�TV�h8����|g��;D��S���`��F�W�NƇ�� Tm3QE�0WC>��������o�9繘/���،3�@x0�Xq�~�G�Y�ԍ����q/jN�Ys��P��=h��p4��p�ui��ǅ�t̖Y7�s��Ϙ����v�[|%���͚&G��o�����H��8����+���ڡ�c3fN�^���2�A2W�����-�r�Ŗ/�[�P��|쟼�iw�:���sYT�4��̪��c��/t���4�Jp2�������h��>km�ط�u�w�V.���e,�_k�����Z�Ζ.]iUk��K{m���eeX��,�h���7|SJ�C{@+���˜&��i�h�z���XXrk�� /�f� ^�L�C!�h���"U��o	�)�����������[|��Y[��u#�5��ⵡ"���~���M,���c��������\Cxa�J���-��y@H�G9n���x��k��V��Q���S�;j�uy�)kQ�g�y�x��!�'�h8͕H)&��-���	��	������ܷQ��%�K�"?��k���~�aW�k��C�A����(���J�͟�_��9{����C���۴�s���P��R��E֞|b�����_���d{׻�<��*��>�9[�d��q	>���c���ZҤI��w]o;n����`?���e��T���k=�~��,؋/,��]�mmw��?�-^	&$��~%K}�c��s�=�Ԣ��E�H��;��/[��ə�8�F_�`��I���|��L ���EI�i��t9ͅk�q	�Pf�d���Ikk-bHQ@�6����; �u��I�S<~[Z��{���=�??�S�9+UVL|��P����!h%��c(���z�}���a1��b���Z�2����\>S�#Ń��`�<��(0h���j�!�>t���H'	������׃�蟗r�M���;͹|=��1�>ڵ|.�h$���ކ��j I¥�3��V*�����ȦOk3��k�J�z�j �,�j�y�X_�Vuu��g̶SO=��i
eOo�֓���������[�\?^�tG~)C��?�Y�/�]�ٙg�n��>�z{�Zo�:[�f��^�Ԋ��X�
�P�����ޛ��]����Yg&$$B"�B�w"�Z��IP����ź�o�׶�����V\��KMX���(UPA@�%����6g2�Y��{?��̓Üs&���f�����[�����7R��n��$���]^���Z��c�5�h��[5�Ź�lX�9G�K(��}�r6i�*�`S�v�J<��^��xnv�h�C��܏�b�'�h��{	E#I��<�T��V��'����u	%�8�ǻ�X�����L� 
�8������	�J��w	͋�8H���w��%�]�KBw北�:�����d%j�c'&�AQ;ʚ�w�}4ǔ�@��Dsƻy"�~Z��0���N���(��yz���������/E-V�� ���Z��S�#ʕ��E֘�%]P	,ٺ�)۸i��ض�JղM��[-�����lp�j+�Zk[���eo}�͞}�U��~�;����l�#s�h�,��_���
��w4�} 6p�Cgۻ��v;䐩V���y���l��uT7������������C��N{�2����>�X�;�0��+�ʿ�Z��7����/���f��6��s�Øwf#+kT$�H��"�A��7����'ϣ�mi�Z�z�84��^�v���6)!$s_����eE+�~��������VA���&ca0�H��#�� ��3h���w���u�ݩԂ�c�'��X�`.8^�ɵu��+s�υ�������<��k=h����]�G�:��?~�;��W ��E3����������G��k\Q�����̄�rX6@�Y�YG�j+W-��+�yC�O2)UISV���u�y��c����`9���o�b�Q���V#�Ϝ>��ŋ_�8G��5�|��Px[3��dj1�ɋ^h/y�mBg���)[�z���w���k���-�-��ڬٳ�����{�M�p���¡B�P�MY}6�e����͆)Φ*��/�C�A�C+��6��ٷN�H�i%[`  ��x�7�V��.��K��I˽����J�����o��d���w���v�W�X�I8�z
���9�o��OE�$�~�Lڲ� e������" �oqss@�#�j�K�wZZ�Z?z�V��-�+Y\�x�Ю��s��Oi���9�_,9^����Z��U�,z�}4�d$���9w�(Ǘʡ�&3��L:G]����Ю&�p+�?������}Bg��c�s#��[��=��mdN����E]d^�r�V�^����,�e˖z1��g�9�y����̎:�y�7���w����Р�}=�}���;7_w�������P���f�/P�=U~�$���KmE���P�3��߱���cƌ�>�^�;���l����YX�~��}CSo?�'�E����rE��B=y>ORK���QYh�W���?���;�/?@��wh�X�y�X��CDE�rs��CWI��i��(��	�h�����|_�?�'n�g��Ϙ��V�Vi쌯Jr<mc%����s��BSS�Ɖ{ro���+��9
�9��^s�8�.�*	X渝e"�wAc幜���I�B�B*��y��Z	�X IK�����Z�\��|βD�O,������pP�J-��0�����)۷\Jh�&�ߘD��.<�T��h<��ݗ_� ؃zn�(� �v�*�%�O�l��vt۔��G`��#��b`����Z5�wt�����?�����B���'��?0�����.���)��w�PŇ�r����7�ѝb+4�����+&tǎmo��lHi�L:M+�� 
 ��[��V�U�`3�~������4�j���b�1�<<?��;�#ԏ���R���� Y���Ȋ xV��h�h� ���(�#\ �����w��g�TbB��8+�������e#K�f���bR�f=��k��}��)u\�1㠕ƈ�!��3��zH*zǆg-	LCƖ�b.9��C(sՐ��J��J� Z�"Ɓ
�D;�7��:4s��o~SO|��P���t�Ӻb�.������{�΂mZ��K��ё��M�b|�?�Z(��1ɦΘi���\���~���m��-�t�I�3����+h��+%G!��Zan�3{�t��"����c��;|/֟<�Q>x���e��X6�	�lGֺ:����R(��u&o�����?��;�Q<;:r������>c��nY��+��ߦ�c�[� kq�c�R����?����d�׿*&�����ʖ,y�^�%v��G|�]w��ݐؼ��ԅ��
��G�v�-A&�q��N���zQ�@�I ��ffa�0
��w�$#�k��.@Ģ&I�Qug ! _�HBR�H��
�8��1�t��3�q��V4Ҿ�}ėJ����:V�q�Xm���i�����T�&����g�4�'Y��	�)T�XT�[IZd�2~܏yc���/��a^G�S�Z;�Gt� n�e/{Y�i$��G�+k��^��C����%!�(%��sϱri��{�~�*���\&� �
��ZMp=��'b��Cմ�>�X�5k���6l�b_��{l�A覰,����#�u�%M���.�>s'kPY��Ε��P�s���<���ʎ:�9^I�=�N�c)�LV���ݕ�L6������ZP?��߮�;#m�IS�~�-�|���>@cp���*Ւ�\+S|q���I���|�	�I� 2|���x�� ��-FE ({Pe��w���� x��&͓{ΊL@!	Iڦ�F5o��`I ڪ������Pb�Ҍ��І%(��c�S<����Yisc��|��u��[���-򪬲H�)�ڌ��=O5c�Y+l|��f�'ƛ����an��5�B�C �@�ɪD�o���܊���=@���*�����P������������[b�u��V�Zi�6oXo}=֑!>�b�r�i4M;r����J[-3ѦϚm��j�j�
�}��k��ǟx�)��4���E	�� ֘񮪃$�]>1/���7�@F@��ɜ����#�������p-p�`��g�Ppq�[\�#O��m�f�*W��w�C�W(��UK���������B���>���F��
�;�x�5��    IDAT�B�g5YV_�R�/���2�/�i(����O�����^;Nk @$������rN㚊��Bi��(0�f/�Ţ�z"��De�*_E�x+��H�q�𾀓|	��POT�~W�6ׁ���2�5`�;C���{_���~�O�u%�>��@	2_rFs,Z�֔@a$��Ɗ��'|�o*�J��7��]&�c����r�s����]-�s��'�Q�xY	����?���=�[�@�M�r���w����趘���Q� �TyЬ<d�V���7[�Be��[��'/��CCUO�*��Us��9G۔��:�wz�_�p�=�d���!l2��.��b�Xrq`�LD�%�}�}�K_r˝r�u�]�E�"u�1��͘8U4y���o���PV^�*�?)��P�A�w�'���#��6�g���)�����=>��t�~ܙ��ģ+ X,�P��j�] ��OX��~��C��Omj 0a�Ӳ��f&���}��"o��3�i�5�U��X%�(�H}b�q�Qy5�V	e���`��,P����Uw82.� ϳbEȼ�;@�s�O}h?5$G� �|��/�k�\�Uc)*l_9|���i�K��&驿��#��
��8w4:�� p��\��^�U~�VI`Mh#�S���3�|�u&ڌ�#a�Ԏ�Q�'ϫPN �P2@|�ִ4����J�h�D��+���s���{,���Ƶ���c�ufҞ�J���~���8 תVM�l03��3�&M>���i�6��_���VZ'J]RZ=r�֚���|<ק?�i{��<�| ;�r.�k��}�<� d�3�Y
R�<d�X��4�D�|N�"~��}),�5�ã|�7B����Y	h���}*�g̼�L�j	��M��W/_$9,���31 VtO�P ���*�aP����������y�Q�i7oݭ�U��I!ڠ]��$L%TR �������� ����DkDp����y>��B&�@����;4Gq�,`��g��:��Q)��V�R܋��Se��K�_���g�]c��͏S#�q
%LT*�;|(�h�|���YT[�8�����P�*��5���fYc�J�MF�h�N\i���M��%��=�X��
�][%z�K�0N�Ԁm��rV�5�V��-����Ւ�,� ����TΪ�iv��ϵ��DK島e�v��k׻�c4�����?�'i1�j���O~�֬Zm���7����~ʂSߟ��1�Þ}}�k��D]ʊE�ↆBX1��I2����#���Jz�|�O�V�̘9��o���_k<�}����,*t.Q�'��	��K8�Ɨ�$c^�b�[ȥ�l�i��f��|i�, �8\����1�i���f�������s��sU�+�CX��N���1����E�v. �'@��@·
R�H��X�*7�3 ,q���� � (Y ��u�w���x
��DК��G ǽEY�V�C�Z�[\9U?U��Z(���������{	��h-1?qKF��|2��sJpKH�* �IDOi}J�ig9�{Qh��yN���i'�`��+C�~��c^�����ͤ�����A���?q�A���i�7m�k���=��S�'YJ�kY	�4Z͟{K@�;DΡ�S���N�(��0'�7��/��/�-Z�w�Y�A�Y򱐕BJ�N��)�(7R�5�T
ڧ���ߊ���-�I��a�g@��ed��ؑ�zh�f�6rp'�����l
�pπ�J5��]K�KE�p��.�f1�%\����z��,�&��k�+-��%
�N�)�x�[	1Q^zY>\[��! >��w�j�tہ��~��k��ߧ6.�)G�@V`�؈;����A|/ �z�
�JK���{�ΕI!�����R�RxX#G=S]�%]��.�x}����x.5�܃:Bg�q�k��r�i������W�N��.Tm�6�τ����߶�`_������K�ӹ �{��+�_�_
��]�� �1g�ׯH;|Z̟�nY�Z�4��A��9m���8vi���@5,�)Cs�j�[p�8O ��	bT �2����F@j�6��9)��'<���:�Mh	���L;�ԤM	|���:|/� ˃��9��:Ց��Ε�(^�Rڹ�M��Oi���j {����3~�����������v�Y����x��4F��"S~[e
�X��Kc+kP�1fXr
�%̹����@V�"��%4W$F����<�-��;�z� %��8�T�Ҁ��l��ֻs�u��CA=�\����;X��G?�&O9�JՊ;|���km��-MYD����h�I�/TJ{Y�1Zl5s��B�+|r��}:L�p�D��ĉ��aǡ�M`(��aއԑ��8���n�&�H�x�w��'�$uК[���~
��EݼM4yi�,8w6���ht6�6��G��1�h�I𝀸t]I,��2��'�]i�a�,:������������g�<���qכ���5��[�RG��(�4 |���d��=�y���%KB�p�rbK�yD`-p ŵ]�I��@?^��;vr{�H��²���Gkݶy�-�ԚC����gX�<d��۰v����p���X�])��C=�ռ~��6��Éذ-�wؿ��ڒ'���	�] ğ�̓�	u�g��-8hC�����+�H{/�S���Byaܓ(�B:���q*������<��7[��}�å��,�$��'��A�%����Z$o0�[�n�|E���<S�x,xb ��'��Sa�X[�5���y��Z��b�ǀ��γ
D���Lև�_����k�1xb�ƛA�I ��0�y&(�_�>�<�1��V�A�q���X�J+�/f5�r
�u� S�R $���� ֕����K1�wAP�+���V������4�����M|�YgZqh����n�`�};]3�=��}�zy�9N��6���6}�LO��oL:\�f�lϱd�j���)�Z�{SV����֘�Ա%1]Sub`!���+K�-�,�$A��l�q�g�U9a�8�����3�N9�6s��I-Z�9ߛ$X���]i��9�L��� TG(:=�|/�1��c��5�H��4�F��X�-Pӂ�~Ah��&-�V`�0��5��Jck|T\_QJ������#M<�}bMZ=~e�s�6z��^��K�Z!v;�hT$�֐Rc��<�^��敟��@9��)jH�C|s���ח/G�+%{:��x���8�=�7e��;�s�\����?�{$��p~���/�L;�&M����t&�͈z�	�{y�x]�oQd�?�B!�!<�)T�$V�4�u�<���%�v2I�"ǖ� �#k���Z�|vu�����g�w���74����h�6�_s3j��OU��i�!Ty��uV��qG��	-�����v�g?,��Q �w�7���s��cmN�/KC�F ��,J 8�2����%bm/�$F2y�1�Ij��D;�D���p��]}-#Y-<���B����I���S��4�=�UP�B0�!k[m	�T�:귣���+��w ��� �t,e/���;�Xo�7$r��wYd�����w�q�\�g�6�Xu�O�g��?����Li7V#}����֑�oϚ/-�U=т��"�R����rŲ��l��e;�Dh��YB��aa7)B̑�]މ1�
e�Uԑs�N�_�ּ�0��lG�[n$l�P��;r!����CuR���X.��a��V~��X�o]�!h�>95����7&o޼s��Shf�8�7*�*��v����,&Q�>ͦ�?����c���wo�Q/�&-J=�x��ħs��?QA�P�֢��(��ck MK�]G�[�}�����^���zҤ�;O�2�}M���K�$�s��]*$��*5�ԛ���n��;���@����_Q�� B���o�ݣ|h������������A�A��AV)돜2K�l~��_y�!�{��_�E�PD��d%��q�����T����	��Z�W��Z�����%�fRV���9��V�f%�}���Ý�MI�0GP�t�J���aI瘮��m��J��+E,Vd�/�r(Um�DҜs�Qv�s����&L���*p�|�
[�jm��9���wtUUh�ߦ�[:������zgʪ��o���E6��s|B���r专�R�y�Q������M�;�(F�W6�w�i_|��� n��f/�,���B���&Y
�}L�H;�ƌ���v�V��"���.��G��o�L�*$H%��]�P7)������J���4�%#� Bat�g"ڧ�;P�3�$��'���_���l"Q���44�v ��ݾ��o{���.��rX�4���_^_G�]w���34a\��^�'����?�����ČG����g����̥qݱ��B���̕j=i����[BC~�u͘q�W��;�8�y�t�|����{����k��ҥ���w��a����;���g��i�r�j�Z�>c�{oY����u����-4������P�L>lj�ܜԩ�_-��n�L�^��/8ߦL�T�����n%�~�͆d-Kel��^��^���1@S�����\k#&�l?��O�/x�oR����ы�Q�)iӇv�&;�H&c�s������Lp��( P.1>�`�w��OL�	���X3���{�񓟺P�v)�E�.�&1�M{!5���a*���E�A} (����J���??h�q�>�nD%��CH�������3n��F�S�r l`U��J(X	���Z�b$���7�#X�?J�����|��|�7����b]q��y���BG�&�\l5ǁ���������e>��H�ճ�/^�:[��'ͣ�"X�V,��Cfx��'�Xj�/�D�\G�	�'	�#����V��Y|�^B6oC��v޼��k_{�M��e�tնm�l+V,�%�?b��l�,����c'�x�}�s���ȍ�SA������/4 �۩�����}����Q��+��K�,�ו���
HY,&z�"@�8P'�W�d%����v�F�l^�W� �>��j�/0�3���[ns�U��w,�Z@���)��wн���)�����[֯��3|G#X��<�ǀ?7E�����}>��	�#�i�A) ���0(�} o�h�����6�( (%� ��J,�������}3YN#�5�w���Oh�.���_�}�dK9����U=|QT�O�-t>���4����VX/eֻ�y��m[69��!3���͵l.o��Xg�{j�*/'�z��?�h���j.��_��?
=�����3h,@*xN��f����J�1}�UJ}�}�f{����򧞰����iV�x��!���?��<{� 6����
C��_�����|�+�G#$=�]W\�<-ş����E��i�b�̵`�7�E�l�V�C�����_��o%)�`���i��Q�	�"�~l�[n���q�u�G���FZjD�#m�����?vFslɆX����G��\�5�wu.c�Ӵ@F ��W�(� ������d^o��G�G�W�.���_K�g���w�!����*Ҁ?��I�0N����D���O+��{���"�u��g�������÷���>�N�G9 ��Cq���g��H^c=#�����g}#�K�?�7�\�Ry�{�a��{�9�Dp��6�?ds�e�}�͞��x�G1��n��P
����9���M�r�8��T_�k���۲��-y�!{��-��zQ|fY�e�lgϠ���q'�j��z8ߗ��e�p��{�s����I�OU@z���	ƥ�H״-�F����"t ��5�q 	��f�NL-5�rů��*���B�i� ɢ�;��{�}�����K.�gD�yN��IS�ZV�,�}�9`�{�+���gV�Z�w~��c���9����p��O'1�D��{����h����5�s��� a��������s�T��5��;�cF��so9|��C���D(?�e8yk�>��p)#�1�ozӛ\������[xXq`��z%k���\���sө�elȖ.{̖=������i塢w��첁����؉'�f��y�z�,�,��f_3���4�����k�N�6Bg>o���]��c��T�h����6uY{�l��^��R�����l��-60h�ik�����y�?&�g?��kq��1� L�/~��&4ϸ�7���dS+$NL� ��9�|�T����88���� ��^롃q$�H�B�����1@?|4e�#�U�(���h	!m��8��m���?��'��GGçp��>����zVǩ���G5�YNz�/s����8��P GB�n lE}iޕ��#Q5�&c�H2��(tX�c��q�OE�R#�۽d��u�gl'5��u��CNH ~rB-L�o��?����������h*X�>�j��p�c@����f������8�k+�z��%��ښU+Bu�rj>7�֮�d�}CV���-o}�<m�<���d?���u!+ 큫����U\�3�����:<�䆯~���O�\�+��_dCfҝ6�_�IJن�v��'{�*@ʅ	_�0A6����*@,�0A�C[ToV6&�P�D���׼�����PWg�h��.\���V[�xbU��u�<1M�E��_�!��K������V���p�bR�$9���x'�h�h���sEg���
e�. �xʿ��}���.��r�_EH�Sf�d�i����u���h����^q�hȝ�P4}r}��a�vCͲu� ��m�\��5s��w|0�l�ga�`�C��/ Jڗ��%�A�p~����ۻ�CgL�I�'چuk�FQ�u��r�f+W��J5c��vۙg�k�{����k�-]��n���m�������T�s��q��?�c��Q�~۸a����;l޼S,�.���Ox�_b�k����m��V�u����l�	��#���&���|����	11�x �-�_����:�JQ�Y� �Z���(K0Q4\0@����<M�@��qBSi`������Y�ȝ�q���]}/��������D�ƅ�u��1�{�IJ������<��T�����d�ǚ�(A���c?.���j�����Bz1�-KNV�֔�Y���؃�����E����$vՂ �4�g�c���aܘ+�p� ��ĺO|���u��,p��"�/���l�#��_��N9�h�1�[�أ60��� |��@��u�u{�uvM�_�q�wM�����ƛlŊUu�����p��3�������o���>Գ�毥v�s�t �Z�V�z�~������n�T�֭_i�}=I�D��-ڪ�i�m�/�`'�r���M6�wh�C>�4z�^ >��?�&'�mTB�LR0L��E�z���d����q8����Z��Z����+�tx>�Ef2���P�lFۇ�G�W)�v`?ҳ ��>�J5ǆ��y���P|�`��)���� 4�틠m)�E�)	7Y��W��9�k�B��6�Iܞ����z�XP�^��i�~��n��KV��^�*[�x��k�c_@���o�i�J��;o���8�>x��Z�<�zz�0 e�=���Ga�v�����~β�N����o�b�r�	Qy}Y����?_ڬCg�'?�1+�,m%��o�h���ݶy�:��� S-c=�A[�j���Y۸��iej��ѫ�O�����L� q��lp���7;��������ϙ��)�ub�w��A|���3�n�k9RZb+��H�w,_zH1�#l�/>#�p|�a��d
)������s�|�|4�ǳ���c�Ɖ^��k�ɇ}�u@���k�|��������5����N��`lEi�]�u�N��'�G��6y�Tۺ�ە�U+V���	l��������w����1k������i�{���}�v�
+��i�N�mg^��v��m��m��ګ_�jN4    IDAT�z��=����N����F��w^�.����)ޜ�"
ɹ���8��e[���L��4g�� J:�xB�	x���?BVj>��Ku�#�>�x�!�G�/*N91����N���������=�C�8�g�b�;��{�#f�Y�kV�p �8���oK�\a����M������ezh���k��j�=����G��V��τN;h��v��U�Cֳc�mߺ��wo�Ri����%ˤ��/tÆͶb�FK�&�;�����~��1�h�$[a
����O,�,e������׻U��H��J�#�x\��}�
b���8rM� I��~��	��磈'ێ�!
��V|SK��n�������ڱ�{L����C�N��X���O�Mq�*CQX(~�;{�R����l˦��ݽ������}#,c]�{G�=��%ֳ��.���6k�l�T�v�O~j?��-����)��%cx�:|���QU�t-ms�εw�������[��=��a+�l�L�f���@����c�©6�9�8@������$ƟJ���DD�"5֮_��f��0��deӡ��H����?�m=~�31�p��V�+ �Xxj�  T(Q�s׭�����G�3!���c�1�X��V�]��ʏ}���O}ʁ���\'J��N�qQ���8�@	�_�q�h�V-�e˞t-ʇ��\�_���`�N:�t�{�)��uX���]��=� \j% �8�VU=�VO6D�,���)S�S����V��k�����k˗=�WS�5a��z�iv�9���鳼�@Ov%�J���D�/Z	�-���� ��N�V����J-s���7�5d�9�q��X�l�+�EV �1�OTq(t��1M�HłA����9���,h��<�x �XޓwW4�"|ؓ���<��x�c#G0>u{� }@��˟gR4?��=^t��T��Ѐ=��v����+�[�J^HH�<a��v�ة���5���<��gw�ү����s`W�lQ�_]��JE��5�bG�������Yg�n�Ҡ�je*؎�[��[��'|�t�T�e;�X���y�ų�0�lU�'��/�ω'���]D�ȩ�yh0,.�>o�1���h�fe�h���]���3kmK����=���TB��b�e��T�#�u���Z!����eK��iU��ݳ����Z�]�I8�	�&��g�P��������,E��	=����ՙ��ނu��ڵ���c��>X3gf�"��t�._f����~ *��Ƚ�g��o��Uw���(�J}��|_����/8ߛ,PB�hRJ�ԩVC��޾�����=U�/����W_�@�ǂ���+}�X����_yHQ
,���ĉ.��9�� �������0�S�-�]�z�gvS���P�b�W�H��0�U-�N۱�k�$B�<���z��р|�cT�	P�ު�p����+��Q��`�<��Hй��P�^������_w�[t,+��~����o�B��G}ܾ���Y���^5�\�~?�����
݅KGN�ҿ1��o�P+�F�&L�I}��W;mCyg>��eaB�l޼ս�j������1hj�v���A$;�ݮ����¦�|���f�����u��E/��pdƺ)Z� r�YH�m���RI�K~��a3C�ocl��Iy�V4��s�єw`̈��Z�ot�kG��hL�	5T�ߎ���l�ќo*9��7~/@�3�UnC�[��O�c��*˺1���F�&�4@�������Y:������<P"�s��@V*�uMԏ*�����^U�U����Ο��:"��G��t\��ڱ`b/S��w��l ��_Ia��vK�N^ټ���!�ε��&{73U�,�"���3"���==Ng��O�������3�?�{U�er�w ��9�|SQv�֊ ��kA�����z�^p�c��G�'�hB=�N \i��$���MD��JU�z�J�1h?�z���ΧV�C���0S%yQ�ᐩ�F��5K�P��| ��H���I-s6�j��o�AJ9��y�X9�v���PVl�Vr�	���v�h�}�{�kK�� 9�5*�9(*I���<�ϕ �2ʄf?�0�}�o��"⪣�KZ�?� ��GQ�\����C�k:�=y�s	�x���8Fu���
#�{���zdN��\=�����I'�uE��1.���}^��н3��gýR�`!��F�w;����߬\����!�������`;�Yw8�� R�l*d䖂êqQ�����'���� e`)���O~�K1P��k0���Ь�Z����uY������/��K<;��z���$�8r��w�'�2��1�uI��nu�������f;��X*!R��#�*!�ZD��9����ƒ{��۝��R�S_'I��:�\IJøގk�{��%PdQ�Y���M}�����E7V�˳���R*����7�(��8�X���r�����%y�w�q��ؒ�] ��v��|�a�8�9����&�KR���_ʹ`���Ă�n��(���;��2�j(՜��10��hh�����©q�aځ%1��W:�����& ,��iQG�k�$��(
M��.����n�4��q-� ����S�3Lnh�^L� %�<cA�CM��%%,Ne3rV	��B*Z�#-���H���i�����4��y󭷸�[%k%�)M��c���;���Jƀ��&�*�;�I<��6�~�r�&�����+n��F��I��=�w�y� �`Zq���)�����gkw�-��땠Z�$9�S���Ny �͟�J��/>88�'�h�=�H߫���Uq,悬b�Q��P'~R������:��4*�uKh'-i�T�d/�I���z�p��`�9t���c����[�a����:|��)�<�n�jA�G�
�t��b4�J�ĭ�r�w&NG/��D�o��w�Q�4p�	��4B)8~B�`�?=}��\RW��O���P�v��1�ƢVm�F�_�E
��@ʂ�7l,0�	��ӤƋ�Ն�����8|���t�Q?5~D[�n���$� -���/�_�\��o�y�V�֧�㿧�6�S\��)�d,��1��3>�C��D���1�ז����+�Hc0�wP䞔Q<�p#t>�񏏘������j�!���ZA$��t�M'�%����.��{/&��?��S4vj��9�ƨ~��0��̹j%r �p��TI���F팉Ŝ��o,s���v�]�a3�q��D#�����y�E���c�G�̹^��_���GE� mC�&	o��%���9|o��mN��;�GμUO�}|���ռ�, 61�<
�y�ERu�&}�1	�?Pn�~ 5�6�Nh !�^c���7���X0�bJ�k��%81VXI��sٝ���c��Z��<vXJ��6�ؖ���5��s-���}ޑ�Wt��>��{����M=���s	����#���[*%��L><Y�h�`����j�P�8(��c�lοE��k����HӚ��L#�j��PfA� �Cㅴεهs�h8��f���3�T�.�A6h�Ī��x�K_��_o��ݛ|���}ڙ�.���K(�H��_�����YG��ӈ7'�}�[�����Z�%�j����p��&��r��`����(��7�_�`ų���ʺֆ\H��Y��]Ig�� σ��:�hr�]�!a˽dep�7��u�[k�v�DϠL�՜�=���/���Z�7���/ņ[�ַ�o�(�MhY�g\v��۽����u|/�E ��Ou���]4
3)ij(q����^�B8y��� �]���B�'��F�g}�}�$�V��6(��������J9h"����kv.�E�*b3O� � Z���j*���U��lp	��h���z�����k�'�3s}@�{�N��h
�-	gv�Ӝ��J�½�������v��L�,��rSI��	-z�	��d�k�	,�m�=�>����
��y�K-�f��ˢE�p����ޚcͫ�|���3��:�_|�cu
E���<�p}���{�ܘ�z�K]KN/�����|
l5�;�m�Gćs��#k(���k� 5�w���5ͳ�}�� �@D�����}���,��U��4r����a�N�c�}��Ĺl	�f���]g�aV��%���ש� Z�j�qԹ,�봇4�X��$���ڔ�`k3K[��N	��G�^���":���7��ɤsP;�m�X̭>��X>ZԊr�i�+C�N��X�m�ϭ1ֳ�����Ƈ�cݐ�G�a�k���W�q>
oe^Y7$���_ �O�'��ց�ќ���F{���H�VS:᮫� �(d�1�K���G���{�ð��OJ�H�5d�"n߮��j�����5(�_ᥚ{Y$z.�����)+V�\:��[�:��0aP�p��q�R���bZi����Z�UfN���ŋ��5�I��z\��n8\(�Z�f3!<m?PA�
�d�<p1o�9d�2�����[2��P|���^��/ ���r���AlA��'`�l�*D��e��iNc`޳��c�T>��9d:k|��~��e����{�U�k:�~K�.��2������C���x:LUX��|��zA�v�/���g�9����E��e#ϥ������+�|߯��u�^X�-���W8�j!J��s�,)*��%�yX#t��3d�Ha�<�Zk�fَP�'��Tj�vM?X��/���l` 亠t��������fQ'�_�iH��gsA{��ET*A���	�삏/�dtuM���m�G�X��Y��5�"r$)����`���18�`k�O����o�������c˪����6
���v�?��ey0/ZC�B(���ؕ@˩����X��<�@D��Ɖ碥���|����xʊ�T8��=��كs�!��}+�_o-�.�ZPb�v�':_�[��["�CG������mw���g�a�C�JV�r�k�o�	C·"ɔ�r�c���OP:�Y�Dw��f�h,;�����eѢ�5��[��2�vH�pS*���<ҙH��#����zz��9��*k��2��7W�?G����i�P���c#$X���A9�c�kԲ��Z��z��3vJL_qSi����3n� V�\4�.n�'�I{$��a��r���D	<	t�ݓ�.}�.�5XG_�����+ϱ>{੓���[N�Ш=|����,���-T I�5�kX�D�L	����eB*�sR��E+A�č�[�#�	в���i5t�#�PX~ �O�?�"��-ʸ��Q
�|H|?�2�}*�O�4�'�@`��P�	��3�-4��#�wIݓ�u���{����I�ä��j����+��+_��L�4w8IY�h�ī��� E P�����P�Z�5H����t�Ӥ{���6w;�2Vڧ�{����힯����^f�45�9"����ii)7ɉx��7�R`�M��m6o�E�p} �� W��}^J�gQ�I4j�l�r���+�%A�t��(����^���{��QC�lҫ@'as׸��e�r{�q�^lq��aD�o��*�u��-<�,�o�%�޵�M�4��e�E�S�vJ���B�ּ�1��=���g̜����{�N^0<�=�Č�8a�k�z��k�>}�o.����pg"���r�
���d3�������S$'}�{�sm�c�S)��G13�Ac�yGF�D��]�����H�c�v�>���>#	����{����Ώ��;�M���T�t~�����Tkgo�"�ⵡȣ|�^AR�	?Q(�$�Y���a,c[n�3��ц+f�|�.�G�A��E����vy8���o�����w� ��h5�/zE��
��=Ĺ�o�g��	����,a���7��N�����3��a0��7�a}�\,��_����w�s�K֟�w����s`g�.���B��f�?���W��Ͽ���/�x|_�I�>�>��p#�-]�G}ԋ�!��X��$/!����!d�&�DkPן��4|�\���`m�FN�QP�u����p�÷Q���tO�c�v�����������d�b�1�lf=�z�{��^=�}��6����@��8�����J���k�j?Q���U��N�8-����9RO��:���^��:�SW(v�c�˾dL��ȇ�ͬX���	����n���d_��?��{�'��"�:�'|ods6y�A�y�6�ݸy�w�A��r��B#���m���5c�R��l޼y6�E^�&��o�f�
Ϛ���O:�4;��6g���2����#���7��<>���C���?����?���Ԑ4 ����E�&QO K��'5�ݱƺ�������C�'-p_ܿ�5�PX+hb�����x�����$�v�s4��2�&`"��}�)?��=V�����}/�Cs�s2Vʒvn��|
�#<�2�I(u��'��4y�Y?��T�z[�:�X�`1P�ΡW�%랂����~�m�C��W�%σ0�3��/���z��1����_�Z;���B����mt��rQ�4�����$�;\��Kig��8��3���[�F�$��Ϝ9�.y��v�)'Y�4h=;�ۃ������>!D��P�{�̙��9�γO<�r���o��v�Oux�I%J���ϸ��`��ٞHu�M7�BQ8� B`o�v��@��g�T�)vp>s���TH�Q����k��ۃ*2{�;�a'�=ޣ[{{lӆ5V跮���xJ�V���� �P7%���s���I���ȭ�
�쩕��uBI �	��s+�K|=���uS�����\P����~����Q�KKz(����g�A4��fO<�����_ن���EG�;����K_�J;�i�����3�����X�Ԟ|Mn5%�I�����=2gh�^���eo~����X�V����Gy �Х,mIĠÎ�ݶs�l�}�)�����d|�_p+�L�^ij�	��B@K 9�@	"\G�9ƪ9�������h����}������ڶ?%�N��J�^�nmw��|���:f|x^�8�qکf����{mӺ56�W0��)�x�\y��@瓊VLuج������X:�a�6o��v�=��ɤRR'��w�e�)���UI/|+�X�m�v����*��d[�s���N���?�K��m��'l��mǎm�ˇ���ض�������/p�'yq����5o ;�������G����f�?!��\Ʈ��]v�	�[�<d��M��a=�M�a#NU���P�6o�j�r�zz����y�{��o��>�
�BCIJ�FS�o���1�X�,�}�����4�i\��7C=�=�Cy��}"��Ya9��Z����[��P�m^�����[6U�t��QT~<�<4)��>ڮ��N�YGk��l�|�mܴվr�W폏>�+�N8ޅ�nr�%j���|�9�9���|��������+}��"��p��|�	�ʨ8�g}=�m���l˖��}�V+���O~�P�f����[�k��v���d�Ϛ�>GJ�C5������1��/�����U���#f٧?�I+ؤ�v����K_�+�ؚ�O�P1�Ϥ����o�W���!�������h�+W�ts�E�v�$oȞ�/QB����x!��(7I�g� P̡j(5���������)��=j
:P$k�}�{��u��V+Z�<`�6���m�,[��UܑN�r�g5�\��8�	�TƊ�)v�Q�ڄ�S,��t���7ڣ�?|4%v�ǘ��2�����g�����'?���wB�����>g���o��(~D"  �t�l���;��C��	9[�f�����~����mɓ+��s�-}r���%�_��I�z��-[���4�.92��`Ⴏw
ok�1�s�e������%۶}������i�t�֮{���{��e�����    IDAT�b�o�������csO8���	��/���o�' Iߑ��kV{$�LH�\�7�����G��J�ߛw���G@�}��Lo�P}6Γ�3��Ph�r;��ӬZ�L�d[֯���sT���x!!���:���9G[��If�[�q�]�MN��5�p��c3�PO%g�X[�k��N�o��o��ˇc��K5�T"�pN�İ[���_���v�I���i�l��%68je��R���\j��D�)XG���G>�e�=�._���ڨh$��f̜��3���7�oo��cY�l�a��UW}�2���Y��������ϰt�h+V>i��`����m���f�&K�'ز�[�O�+�����p�0���D�Ш�Xl��p-8@��r ���`e	s��8���z����N�V�K�z����1���Ͼ`ݣ��š�rѶ�_i;�n�|�h��̥�g=�W�x�������?�c�z�6a�:�_����ǖZ&��������/'� ]�^�erxN�{��]����T��}��\�(�|���=���7?��O?ΦM;Ȟ\����RC�\IY���Ǘ��J��ne�Q���������W��ei�z��
0�q�o���P��c���|�*������n��[���e��N��i�2����W�uk�8�j�v;�Գ|1�0�pH�R"���p�͋�uHn�{��_zM� ��Xi	q�X7����f�����5(�u�����1߯��S-�\�߲v���������<�����pNJ����MʩSژ�+�.;�����I9�a�6�{�I�>{����w)ɐDټ�U��K/y}=�����Ɗ'�+�6��|���n�Gp�Z��~����I'e3���_,FLeϜ��Wm����M�ի��f���_J���E��v�?s���,^����1hޅdls��9�=퓵��{���Gl�d��J���l��2��l����D��Sy��9`�W������ۼ�^��=1�E�VOU�X�Q���5k��0��;��]w��G�@ H�h�1~�����2�u����kd��x&�M[�0k^e���f���_.Yy��6�[e��[-�*:���s�?r��-D�0\2m�s��	��t6���W��	���h5�8zF���ڹ��m��]ٓƯ��4���>X���Ϗ|�#^�{�f{�ޟ�ԩ6m�[�&��j�O����-yb��Kۺ��N9�l{�%o�l��Ճ[�n��>�4���E��,DԠA��Mo�y�βJy�V>��OD��MV*S�+0qZ���wز�k�З���>��?�~*�+�-�_ř ~������淿e+V�p�W�Iu}�Q$������ZV�B��~�8�$�U�V�+ئ묷��&�3��]��fB�$J?�Pޡ��Z13�fqdh&di���o�����%K<)ʅ_�#@�Q(�(�W�J�ñ?�[��Ź������bG�9m5��F���gj�fգֻs����PiЊ��z��T���A{b�S�}G�]~����G[�����.[t�b����w8���uj��L�,X�B��n,��90�9�ܳ��^�5��|�=����z�2��-���UB�g&�����)���'�EA��?��?{B��_u>N?�tC`Q@��G> I:J�V���D�rm�6>��`��M��@M���ζro��};mݺ5�ӽ���L(�P){�j)�����[��pJ�lαϵ�3�r�fk׬�k���_�[�t���bv�m��b��GV/����|x��.��"O�BK��Q��i��fW\q���u[G�h+�z���1��3��8M^x���6ڑGg��=զr�z������
�Й�f+���)��Ќ�'kNN �-o~��ܼi��rY{쑇��?�gO=�ܵ
�M�2ɘ�SO9�;�X�0�5��~����U�a��kQ��E/z�O>���'�}�l��yZr�&ܳrW�?���bT�=���-��sfϱt��e��n�s��8��R&�v�5ۤ�����̆�;x�t���ٯ}��v����Kg3^<n,���Rv�BV�s�ᇻ�O�{��6n��A������ܕ<W�pL)���~�I��mp�����>۰a��{P�3���Km�aG��I[:�����{��7%� ���?}��?? ��/X�`qw���f௸{�e�v�An��>���b�y�F۸q�k�8c �9�g۔��Z���Jռ�%}�"����,t9�X8,~QM��n�A	 -�����Q���C�G`�G@>	��؇h��K�������i���JRO�`;��7�{�dC� ��syotB��2Q.y,�P^Y �[��f/��#�K}�TЯ�kO��
@�Wƾ�J���[.���'٤�]6��ok֭��[6Y�@�G;utu�o����������sg��46l�d]��R�|���h�\CA&�:�d�⬁�g�,jF�Y���-W�w�������ކ��rI�Z�B�������� �-��1�ݻǘ3~�d�� �>�F8�N�T��x~��E���?OS~� ���b3�\����/��k륤�m��nr�q��#y@�=��I�1��:�����_o(٠�`a�D!,:)�X�0V8f����^!����S�W��6�Z�����Qb�4y�$��N=��<�v&v��8�H�K9�t���v�]��D-R�	��#mGf��'���\n��Vw��!��}����kk����
�=K���c���n��ִ�Ls]V��U-nըf.O�2��}��| ��<��$d�f|o��q�!��)��B�k���.�GA��=��c}c��@_g�	�N������>˻{�96i�D�˱��W�xwa�=��?�w�����������颜�E��¥M����E��rJ=`�Qga@�I'�d�6+D��.e�n�:{rٓ�uTke?��^����|���������Iǜ�$���/}�^�{�g�������Ox�F�9�:�Gh݇it�x6g>��TÊgv�(�\:X��%}�^a�����pކ���z�*�M��aһ���b�Ja�h�T椌QK�ݶ���H��[n���<x(�SԮe��1Ӟw�q�QC���ֺ����I��� ��Z2��g����i��l���-�wh�B�K,��*�)$ӏl���W�&Y�.���+�K�I}�At!�$�aʱxT/����Z�*?�7���l���z��T���(?�o�G���V�F:sU)��M��Ϯ�<�(����@��Thv��tٓ���t���l�T�Mq�q����.��K�ѽ���5�y�G��H>�},���>V�s�\.o�	���A�� 4h3h����i�jq����=P��Z:|ہԮK��z�g6U�V�d�0� h�w�����/�ܣ}p�7 �_i�m��6����ydA�:_�$��03�}g��3�v���iQw��=I�zvvҌCᇲ�d;�c��c͓�"q"���n~������s�]H ����[�s��J�(t����9��\�<��Q�~���Iڵ��8nMg��Ww�ۃ P���H����8�"N<k��W�pfL��������t�v+��N�'�^h�� ��&�|�6�I�Rr����gqxƐ���
�5{�Z� ���\(t_Ҍ�i�hw�4�H�HׂD�F8�QC&#�i�${�(Xh�p��?�� Q�8mt9��=��,�F�R`���H��I{�������ꫪY9�Te3N}%�qR��"����ZXm ��3�;�Y�A�|b*�N4�D(Ś����8b%^+í��÷��0�`�?���`j�T�H��r+�|>�A3ޟ���1���F��q���u�b�|��i�E���@0r�E�m$�4�a]�8Gxb�oT6C�]��� ���[
݅�5�Ȭ�al0����ݵ�P�C��&l܀lB�b��y� H�ูs��_����G� ��|����ځ7k'��c�s4�����"��H���6����|�p�5J���F4��Q	u��Fo��s.s&
A׌��Aɛ	��g���]@0))�b ` 2����
�9K~�z�9=����]�曗@������/З(��I�S�%
�5��`sW���� ܓ�I�fb	Z=�����@���v�q�Ջ�)��y���k��U[�8�!�����hB� ��ڰ�$4^��a��*��:̀?~�x�Ŗ � ����b���;��š�qmX����M.����7��4���f�Цiw��o�}sd��j�Q������
i�~�H#��$:�g?��Gy��G�^"�D�i�wը?잼a;���w���e/�g!_I��Hӗ��"�#����<)%Nt�~��H���zaTJ��y�4�yXL�7n��S)XJ�ЇW�SFN-�^EK�okĺ�?�,�?��<h)��g�����������w A�5�@2v�{�����o���/�0��X��'�ä�$d��7"rX�h�Тb��Do5�rI�m#!�nc����O�n�d~�k��'y�]v��#�S����6��V~g�5�׽��노诊3��)ϭ�h�Q	�=��9</�Bx
��1S?��K.q ��C�(nY<�֦�T�?�C���~�v�d����� �IɆ䨘�ј��\���`l�I�fi��.�b�^`� Ƣpȕ�В5m�����beLc������0eLe0�g��Ɋњt��,��c�. | �u���8�9o�[���mh�с�������<�MT&�DX�p�C�x���x�Bk�)�����8�+�h�l��*i�!��NDD&�z�}����uɌ���{�J���ҾΫ��"(ش*�G�Y1���ַz��O��]�W`�����2�5XK��r������}�c@V)���F��H0��#Ǣ4} ��������=w�W�����Dah/����� �m;��Ԧ������O��ݿ�m�C��<�( ͵�K��i`}�=��z���X��t`�f�i$�W)_	�0t)��`ķ���8��bǵs����G��kk��%��1	!�D��eq�~� �`���h	���e4�M8���&�o|�;��m5L��Ip�o��q��(�y��۳�c�����$+�ͩ�
�CV�Ýު��/j.Q�Ma�d�V8����g+A�O������$�(,Z
�9Gq墴(6ȹ|�(�z�?���τE�j�b��-�,}�CH'�a�/8�����]�v��X�$�R�4��ź��[5�J2�+��#h_+Z,�V1��E�P�%��1pBkС=�C�sW�u'n�^
�<��$�HB���{��>M�R���Q�X�������^�W,�i����6|aW*aMS-����r�4�7���A,�4��c�\s�5u��V-$�<�?��@S���Vϱ��٘�?�,�GqB�G�d��%4��[h�1u�9n��G�ٷ�v�����_����Ų t�	�(�9�:�/�_>Ɓ�~��փ�����pD����빗Ʈ�4���@K��%��"��=�&9!�z�g���0Q���[o[;	����FzW������*9���`Q��^ba*�w�Iiq�I��	��  ��
H�s�o8����U��g��[-�z�q�V^�_�G1!Lrp&��X,{�	���PC��s��`��g��!�h��ڀ7�i;N]����5r˼����'��x�R��OPS����$υ���UO9���M�vϾ���%�{wzI]4���6&sR.���&��8i�Gċ4�Gy�#4H�{����2̳��4ƌ=��C��/}���������;�0w6�p�����w(,E��x��~|��O���1�� bE��p8�'��P@x'~g=b!���3���|���e;�Ph���)�(;�	�q$�F�_L�2�ڇ��~��J��E�J�c�j�;�9�5�����go����6���˓!\�s"Z����!<�����۔t&Ҋ�r�'"FJ�PցZ>C�%Ky"FH� ���&�����L�R�Y4L;͢FHk�f�x�21�)���SO�%�i���������/: �>�E�
`����6I�wؗߏ�1���	E�0?�6m�wN�]xw
�Q�	�j ��Z][��\@IQG
���s����������w��T<�a�5G=V���U�6�d<��z?E��"��(�����d��iR���Md��L�X 9���=���Xʖnų�7�F�  �<Y�R��(Q��bv}�Iu�l�f�:��BL���'����o�g�e�j5/���nj|@��k.�vO��&-.��Ҩj� ɏ�3�K1�9&d�i;�?�6W� k�5��/X
C#BD=V�XQ)--J�G~i.֕�;@qJh���Q@��&����m���x��Jh|d%p<�+�z#��kd�����w�6w��	�JCܟ�'���?��d]�����|�󰁪0K�ħA�1Q��X�_@��KE1�5[�����+SV�q�s�����$�+P��8���z&t�_U69�DU�a�Y��,+1�z6����`A��C(���<�1Yj��O��u��'�d�7���}VhKz����P�֮]��@��t��%���'�����5��o
=�5���i	�_u���PaS)��c�����;;;|a �;�&�@ ��O}�S����|w���b�V%�BT�P�0єp��PBVB+�'II���Ɛ��p*�P���'@�;�/Ĵ�H���Q��9�Je�����@,����yVE^�&y6Y~Ҋc�E`]�I4W��8=UW�x����@�gx뾚�v�'ZNjY�. �!�MTǒ3��;�·R�>����{��)Q]�J�:���	?D{��V,���yq�c˹����c�'�k^=�GN=h�K�^��z>�jmE��AQ!/��$�9�Ƹ؆�@�?p{�.\��B����?]S���>�>t�,��9ȗJ�t*�<hK��o����cB1�f�~�kV,g-�MIF/�a����;�vXDT�r�Lf���|:�쳝n�)�8	�j����P)8Y耇��:�
�m�}�}+���%s�<� R�x%�(>����Gs]=�"������tc���6lp��:{�E+��*���=���q'�^�0)p�gfM���;�Qk�[`C�a�H���`1T��o�����$��������;�$K
��X��O�AEO|K��z�~����y�B�}	ʕ�=���x��9a�u��N���s����~��۶�p��k���7
=�l��Z�ڏ9�h���WY��édS�`۶l�%K���֯[W�+���	�og�=Ϟs�qf�഑FF	g&P ?^��� ��b�U&??L_��|��\�S%P��]W��fϱ*���<�Ѱ1���}wa�h��� پ8���Kt�������AQ�SY2�c-V���~��� �.�v7cރ�NxQ]{��㋢Ě�'A���)�/F��ͧ?��\P��}R�.�)'i;�G�]T�:��3�K�����T�Q�W��(�/�fmA�~������;v�w�̛7�#���k/��^z���O^lV�X&]�'�\b�V���Զwo��`����{��v�igء�fCŲA��w�u���e���.���Pxw3�VC�c�:ʮ|߻�R�l�҂%[�~����{<�'�	�#^,��P���*6�������rV�~�eJ��� Ŏ?�|(�a���.�Q���h�8�����Ƅ;��,�����Ak��׿�NQ�nc��o��h�_c�@��;�ck�x�V�_�-�-V������>h�$�)}op�Ҁ�����:'%p@\8��'�Ē��西�ۿUVk���4x9dꣵ�e��4*ψ����x�b����ݲ�#��+�^�w�(B����A䟀�j��Wi s��W;ː��l������ۭT���N�J�N����vX��������3gz�2�/}�Z�0��8�7�\�](�yS�'ڬ�=�������:�+���G�\�f[6��m۶��Ѐ���&��d�;z�ڂd    IDAT��3`���]����ɇ�����!M�@&��w��Zil���\��_���9�D�Q�5
�=tl� #4�$q���}Ќ�Iʂ�F�_ ���}����[�h7���z?�񖦪��
9m�c�pH8�.ມ}�M�7�_�'
��E�ٗ���z�s;p��g��1s�L����.�3}b_M;k�s��wQ/�۟�2�4j|"������]���wgw�}�7jU*�? �/�B(�.������3U+�6ԷնlXc+V.��[^�D��l6o����y�����\iO��x?�������:���]��bw���f�_K��G�9�>�����@�M����n��.��� ֮Ya۷o�\��:�]�u�[�n�Y���o��N8Ů��
7�]�Z _� my�ƍ��H�yի^� �{*zB��g����*}��z�ȗ�ǚd��T_ ��
�����w6 �Ɔ��;���X�o��}H����w�+�BY�� T�h��rG]+����D�z�Nq��G?�dAU�P�E��u��FT�	�ڇ��Z��������o�AH�r=�&��g��%�g̘�5���|ͺ#T�dAA��X8c)��	��ՙ�O-�AC#�3FPP#3���07�&NX4&�q����d"b"Q.	J�F�^�`��@7�s1�xM��#q�Q�iA��޻����WOq(��k�jY���t�W_���<��>�rP�x�Y��M�Jc�����׭5~�ayy�ik��wW�o�˫͇��7�1�w�W�A���u�Ŏ-M(�i��H���<d��u�d���_�5eʯb��݂?�燆�������M7�p�|���<������Gc�MC�G��9f7L4Ti6|LPg�Ix�f����QGO�- ?�E����8Ё�<�P54 {��G��ի�Xx��J��^fF
�;�?��?}�o���Z~����[���Y�%��:�d�fu䘳>p���� T�8w�~0J.@�9h"�S���"X�6�M�EO�%
ȋ�"@1q���yꩧl �@u��$��3 ��/�Iu<=�("��RC����0�a'ث.��0����7W��>5f}çf�A�������~����ֽo�����bQ[�ߚ:��-��K��<�Lq���/2ш1�]e�������cL<�l>��cӴe�Ow�+LӖ6��ǟ����yo�f3��/��.���0l*�@J����ۇKI:"`y��[-=|�p3c������8���,m�S���R�A�C�台�.����JM7�dG���k]�G����g&���M�TI!�"�'��-�.�5� _un��<
q�|�X�d���Y� �|����_wQ>�f+�y�ր{��,��^ u��M56����9r�5 �V���QG�6���}�|P�.�$a�zM�ii��-M���%n~>w����kk���^�j���g[�IS&��m�$�����u�Af楗������d=�����<�$����47��`h(j�������ΐ���Ō8� ��N��\s�]t4�ܹs-/�;L�>�Eê��&��c�)�:@P����\௳ v�
�l�����MK��ϢH*��1��m%�FA�����V����hH��	2�~�Q�Z]Z��a�����~��t���C�˳᧒8�X��2y�9�G���;{Z�s4�C��|��]��3G�=���>f�wM{'����6�xȼ������N�HF̜��7Ѳ*Ӵ��zZ�Ye�?��UԖ��)S��/��P���G�0�~t�ikm6}*#�ŏ��i���f��LssS�(��ټ��ԯ�Ĵ�yf]}�w�?��*�}p�(��h��1cl��,����F�0dlD5�Rj�
Tz�i�/ �2�0Ȳ
��eec�0d|�,l
�y���}7�ߵ����Oh��;��Ϻ�R1�}�]̅hy�<X�Z��]@6S�Em�C`��N��@_���&�y�1��c�W��۾� ����Ƽ��-�67��_z�x�P3`@�z�*�mNUl�������۫L$��l�3�c�8�_L�>5�ݕ������?>h��/Z�����s�zZΟl�2���!f�W�f�;oϴ����+�j'�j~Sf������6��Έ9���e��T�e~'�kN�'5��xW�/]��*e(��\bU"��r��)p.���
��B�jN=�T�{饗� ����L�w�cU�?�%��^��N�F���_)��.\h���gk���m�R5�Kɳu��s���=7���+��Wz-s��o��k;v��������%ւR�<���iv��u��0��m:y[{��:&u6���'����]mZ[�滧�iFr����k���^��C�t�a�Ǉ|Amm�}E���LY�5����������ϛ��C�d�;[�����7�3ﾻ�������ܞ����io��ƦN3쀃�q�Oܦ/��Y��<��ݨT2rF���*
c��	E--�=��rnfDO�?�������W���(��{l�Z��(�02
�10 #
��5R�]�$'I����V ��G�=���v?`��;Nl���nO�
	��||,g/�g���b��b?ślX��Gٲ�Q�jAk
2���V�����u+͇~`�;�MUE�54�imQ��xɈY���f���jL��l�����y����r����Wjݱ�/Z�h�=���'?�;3�Ӷ��:�/�O7t�����g>��`ֽ�����?���z��N�
E��Qc̸/kF|�M�b��T����c�*Iכ�'k%�e �/!S��Z�͛2�}��kv����g`������m����ݢ�l��a�_Q�����R��B�?�F~?Z.�>���2(���X��(Y�
����qXQo��,�G��œ��>���Q����I��)�FԨj3x�D���7&�n�Z���_�����^5��wXs��:ZU��|��c��8ҔU��:���j���{MWW�Z���2h�E���w#�?�;=��O"x�3<�\p�~��6SQI5/�.v���&[�a��>��4π�M(L�0����8}6���S�G)�Hq#�p�|�@_���������y���!�s��P�}uV��J�T���ϗk����@���J�
HRTUc^�o	��S��8ܞ��M��U6�/�`S�|jW@}��/��v����Z,0�o2�ԟ����~ �?cٝW�-�L�K��U� P*R�M`�ޢ�T$�B55�S���Y�<� ˥I�$ݓ�l�w�3��N22��0~"}er��*󅹄��ء�m�Y�V�N���$9=�Z!�x��}��+�@�t��d��P晲s�ռ��u��4�4���I���|����oжй7�p�Ut�r�<yW�T�Ϝ��Czx�J:��x|���wW���B!�|�!>������U���o[ϊq�zy��4x��ŋ�Ut�����EA�Sy����T��iXm~��L�l(����k�͙��A8�� nZҲxO?���JQlmb��ֳ��ci۾(�d� o] +��o�l�w�y�n82����¸d�Ӧ�	 �߷��4�8Nm>�	��N�� �%����Lj��	��1Gw��{��ލ��� ��\�YʖM+�W��������)���.��gP(l�p�m�ؼiQ��ś3^��s�̖R��e� �|�?���i�(i�.G
�"< [�3�Ea�1�ָ [���@V�1'F�t�_����A��}��-��J�=�5/R��Q�F�8cE��9��T�=k��>�2{Q���x����I��}��r�`/
��!7_2�Z�Ƚ�KH'�I	�=��y�P��u��9)e>�{)л��@3n�eW���d{y^29dА鵵�w�O�2��Xl�iYi���^r�%i�P���2�u��p�b&GY�dA�B#+��E>���m M�g!N���D�p_���{�9��]ֆ�g����V��:�'VY���o��;����,O&���%o�k��l[��WXA����[o5����=�@�a	o��
�@���)�٤,X'Z:c�1mf��OA-Oϥ6���U�/`�����R����n�=2!0���f������<�J����?� �?�ܒ��u?���+��s<2���;��sm!# i��3�5���� BN~5�����IgO������H����)����d�k�0�k���y�f���4L�N�b-�Ħlz~�Y޶�8�:s�J�3g���@>���yF}�����K?��/�j`
Ɣ��xd���<�U��~;>�	�i��HnZ�<d����u�.>�8��b����2�m(ֵ�N�,~iu*��,"`ON?�}�m,hr�9T�ŕe�=%�,�[\"�c��h6n1�Bl*�q��������m2��ҳO�4�o斲�mO��
�;u
����S�>m��WUT����y��l&)-�k���x��h���r�=�	�]*�g����q����7�^��\��Qq��ѥ�v�`�x��z�H�\����SbN @��w_R�Re�} 2d�,�=�.�(�~���chqrޙg��>7Z�>K\�b�-�1�Ϥ�d���[6����c2��s�O��g��{}{�F)ɪ�QCCq*#@ԩ�J~b����w�� pƃGKJ7��Fź�]�}������C�e
Ƙ3)>�xP d��ٯ(�[/Y���d�Ew�O��(��N6�P��&�_ZWՋ�����4��>�$��92a ���
S�xJ���j�An�� (
E�k�IG�*j�T	cM ���u���J�rS0ڂN"nA�GQ����d|x"<'9�|�R۸�@UHV��R�6������*�Y��&��
�G�bL��8����]�Ck!��뤸v%��'�LjL�����di�&s�����҆��|����7�W<+� ���E7OR}�1�wJpd� �6m���3-��d	���'�p���/Y�ʣWF�֒�g�jf(�M��?8��,���3�z�V�T�2�}O��`��KT{�q�x�������^a_��`�^c�6U��Ŀ�E�fƈh_�oK��simm����)S�b��og�d�Xx-� �u�]Nյ�e�sf�YH�G��ʱT����D\�xg�ϱ�\���?��u��a{k��`|?���|��M���?�����pc��bG/rL���	@]�������������B���y�~ �>�:[�L���}{��~}}�H
R���񂠜Di���������"�2t�;�ȋ���Yw����nv����3�N��q���F@F�*��z(}_YW�||�Z��|?^�&t�,X))�����:�w��7X�^s�g��W�j�	䛗xz�${�1��Dɸq %> ��)) "�^Jo������/E��3�%Ydb�0�k֬�^s X�c.�,���7M5)�[ލp@^�"�H{^�\�EJ�>��-�������ű��)��_���@�)��N.g,�ׂi)3A��I�
�[�wJ�k�
tt��o}%ҁ%��r�c9� �Ud,���J�g��R XԎ��x|��tM�����/ZŢ͐���O���>���
��e�5�@���f���l�o���<3|�a�2���gPX��Z�?�Q��8k���ڂ�9����z�QGٸ��5�*��}tϋ҆:ԚBy�(AY��R�2p�K � |�M��K<��ISK����r�
�?�D�7�H�~�<���=��+�����9k��e}\�'��ε��KE�6��c��갺y�|])��xc�l<�ﴷ��(�[�F:��N����b���g~?����Am?s���a�R4�.nHaK!
oDm2���d e�=�Sy�:s�E�*>�2��X�qj6�( ��L����ܝ8�dIZ,�A��U�h)��7�{��J��od�5�CX ���{ �@��թB.m�*�Y?�ļ���nu8d�w6��!!�6c�!��象� �x"����������,}ι��=����$_���e+�U��`3纲A�lN?�ck�[��c���UJ������������V��D� J�C �~D��PV�A�+D`��3Go�����!N|S�f��D��p�}Cn>�$0��(*�/Y�X��/Xʌ᪟α�*'����d��k��"� ���������s.M+c�k�RgϞ�ND`O�	�-ݚ��d^dy���Y9��h<cP���衇ڸ�G���R%�̢.?�Y���\cEϡl#)���Z���amm�m%�O�����d�?�kd �X��d[ @���� ��ȹ��z:��H�:�`�m(��Q�6֩
L ��+Ț�Z6�F��~b���2b�� d_�m�@�����o�_)����Y	xc��I ������Y�� .:��� i��Rb�����X۠5b�?�я�gB�(
O)�xU�.2$\�����s�A@A2_o��Ft\����͂s<����{sv4��1��O ���� ��/À7��IW՜s��f���|�i^ޡ�͟k�H�C�"�,zf�����]��+Gm�0�JBI
�ˀ�U2��}��naݭ%����_�?V,��SD����
�m�`
�@�2��7����s�)w�7%%e��r�-�2"�!P�����L�����Oa�����?c����k���8�kg���O�1,�Q�F���41"����ǈ@�g��W2�I���\?�D�Ld��Vy�J]���|3>y��_��k�I]�O�N�VLbW���<��kkko):�<e�c�����h�]�0;���Y�JU�u8F\m7G�;�*�{e)�9e��9l�N2��;�;,�s@�Ԁ:Ԅ�����[+?�����9Wm���l��--�������Y��?��mV�G����W�})�".!�������H$}�D�'N�'�W���qO�X�7_�����}�`�h���В{����ߕG)�P�W4����7{��1�}�����̪[�h^с����o�&���O6�w�'PKJ��q�A����L�/ik��A�?�?����4���	 �^�������F��ˣ�>�\q���anPrk 7���	����s 	����K\5��B�?�r.�$�W@� .� �,(�ݦ8�b>�d�'{�TfёPrx-J��	�fƸ�3;�������\�����(�Cr,��Y`C�� ��|Emm��%���h,#,������
*+�$|�ff�*���m"~�}6ΟTO����(`� �7�'=��C���( ���PN��p}��e��{���x��,��Iٜ�����?�NcA2�|i��Q`�!��CB�3$艵��@�9c ނ|)��A�}��'�M�m(EdIVv�\��v�.���)��w.�_��x�����(h+�'S��d���Ʒ�ͮ[TwS�P��g��ם���5bQ��[���& ˆ<���m��
oد���dc 초����-��!(�!Ç��j��T;2������g�W|�8X�>A�6�_�	�����	Z�fX��z
w&�KcA�'���R�$�
���^
��"�f��W�&�C��^�_5��,�w7#&׶앩���Q�x��񳁿��w����*~W��(�ނ����S&�6�b�?�>�( ��<k,,�P�Kr	�6�r�*/I%�|h@��*<�N�Y4�8)u�M��1��M)\+�%��_�J������@�o	�}P͕��Z��1!�MX���?��r}֚���Ɂ�'�/y�Q�ɋ葇ӅK�c�C�4oi��#d�'�T�jŐK��ݲ�1n�I�t-�\��˂��*�E��mo�zO�[��?)��CO'qw��;�_�� �y��6���m�6�v���KdEʢ=��al����w��%ݓ� R���,.�
K���'e����w�%�{˟N<�B�?�?���rD$�Z6`���`i�    IDAT\j�'���@J������@ܢC��1��P.j{�ߩ ���s�1��d\1 ��y�.��<���������ɤx��D9�j�He��.R�ʣ���Ӥ��Naw��z"�-j���w�9��������:X�8�^X�p��9V/	�@��ķ�M��|�K/1���;����{��M/��\�2>�_U��L����](	��9�\h���� ���-rÒ�(K=d ���v��W^wwy�=ɔ���{s����3�.�e���R��t% ����yE:F$��y���/���x��������Yg���/�˳�7z�@^:�2���q�SEn�<�WM�,�'�|�ƕtɹ
����E�6��M�8hGɂ����ރ�Ҹ�]�]�y:�2��E�a���)Si�5��
�_@Z՗�'mjDux�(�Bȱ�iŠ�Mq��բ@-�y^ �9�?�n @W]lF5�S/��x�0��òǺc,�r+���/@�kh� �����k��w�A�(z������]EQ��/pI�d�駯yU]�LGb.s�*	? �,B㩫+S��52R
�x�z�W��ǖ&t[0p=�} i��B�P(�G� �T�r����}������9�w�F��Y�ъ�zRT�5j�o�(V�+<���0��������ŗ�?iꔇb����S�?̓��`�=A���b8u�+��T� -B(���-��O��=��-<?����<��s����K��d�;�?@��/}Ɏ�!��q�3�=\P��ML�7���;�$�K��d{�m�l3CRV?���~�^
@�� ��?�{���ώ�K�S�bs.P�okB�/T~r�F��5u���]d/�~��;�3�?��24ħ�� �mj��R.R&:�:�X{C�=�<��C:]L��n :��>�߿�GO=�D�w�<e��i�5�!��)��V:�
P#����\RH���XHV���Xx+V�H��U.����	����`s2ר���sp�ƹV�I�5���a�A?���h�"[�K��P��#&o;�KV��)���y��S#�<��؊����c�  (�����l�[)��v�gw����u+b}�I����#�ܐMƩy��� pU��|'ʜ@$4�:X� ��c� �(2��3BYI�!P=('��w����'�H�v,͚�{f���O8�������ŏ_?��S���5�Â��v-��@3�� K)�XH_��K��B��*vt�M��f`#�7���j�q�]�p �i)�����e~^�� Y]�8��a�Gi�P3:>�s��w[AwG��T�BQ���Z���P�� �m%�_�M���m1^x�U��T��ۄK�/V�w���a�J�����j�u��\�C����:~�Oz����O�|�^ �뮻μ����j��?��F���;ڲ��i�9�5�a�o�
���{�N�U����S���"�V9D�v���1"`|]��;����g^�0����|�]����O�')�vO��Y���*�d#�	A�{6  Ϧ@�-�ʝW{�̞��VIc.h"��s�Il:�uF0o���ҍ�Ld|6^p�9���`vu���#��5bx'��k�eA��I!�݄�/��T��\p�����r� P���S
�>�\|�V�*O9h� ����i���h g.�I�k�	�gm����?�Mx�4�|��Nu�d�-|��U�(/Q�Ɍb���.����j�����l=����x�s��a>�У�)B�r[cc�=�~XX�x(����mm����aWf�,���7��T<�VV�{������8�b���ӛU�� ���X��lB62uӗꇱ1F�1��6�!���(*p��#�1�?���R��ݼ��<��)N�˟��g�.���,D�e<sQ�r��$)�C�s���{�N�H .OS�G� �oϝG�U���2��N[)-Q4���߅|�{d\j�#ߜ ����I���]9�U.�x�u���u���o\��-���L�n��ƫ�T�OgJD�v#!�X�X�:��M�S>����tK7��0!��'���@�?�B}�y��C۸��5�Rg�jL��;����+} �j����Ac�Z�j�Z�|k8���-�K��6P1�?����0?�?��%�-M����8�Y2&o��e��d��1l|��	��t�WkKO(*�m�>�g�)��ؖ�Ke~rO�_^��+Y��TRyԒa�0�H���>���[����4�/N�k��������oO���'�3m~��!�m����K��4�":(�'V��$]�]s�VѲ�]�K�#��Apw�M��`���i� ��z��d��]#���Wq�֦n��.�W'11�dz�y��f,�yF2MHC$3��J|�Q�TO8��LJ�J�eZ�C�馛�x�����9Y��b1�7�с�2����x~h}WZv�er�g�X�(`e6�5�<gbܬ��;���^����w���a��3>,h�V�#{���O�~���z477x�7�y�O��7��Ͽ���^_������W���Now�Vs���Pv9V�<��5�  ��'A`0��O�P��݁��YY��=�!��( �� :�Qx(�8������K'�i��o(�e��pjn~
��W�=�%����g��y���`���yꮲ�>��������ᕒ�C\�s�Y���1�8Lf�ܹ�������J����&g��w�1�ͳ�<�[�w�ڢ��|�G|������l����=��]s�����ٰ�e���8d�����)k$},A>� �H��f\46Sa�t��`�ɂE�͘1���~hSr�� ]�E�qh�[Z2�0�^,h�rt=�B �����O�Q����k��?���y�I�ĲG��ƿ�� �W���Jnh��}d��k�i�X�6��mW�|D%�g�d˟uW�+��θ
����e7Ͻi�	�����9��˗G������۾� ��"���D覻;�+�(>�wQ�*+Y@'�7����lyv���H�� �A"*�`����)� ���;��������aEqo
��P��>H�$�"CF']1&�
�����߰�I���u�.�ÒgO�g.)�c�PH�A� J���w������$���o[o�އ�=�3c`Ȏ��x����.Yzaw���3��(��O�x����Y��P�]*�W��-vw�����С�d`(8���Im(�_�)$��͟6	��un��RN����c����= +�-���q= �L��Y�����KA�����Һ@ֿ{���f���8ԅ�o>�Y�FoZy�V�?��5'�S�H����'D�
�WZ�^$��?xg0g�l��T�2��ֶ�	��y��=[���5׌[��s�Ps�ҽ2b�Ӽk����_i�n_ײW���b�\|�S�gf]�gm<�,�Ϳ��J������a�Pm�p�B[��D�?ܿ2F\�E�|ƯϺq(� �5k�=xE�\�	TP,��]/��C� ߮'�{*� F��d�`TA��8���6̤%sp
��<M� 
��ۓ�}���7��Omʭd��.���rS�Y����7/�q�)�?㌕E�<��c�}��~S�J@���}������XG��4Qt�jS��|�3��<7cb������%�����8M�Hl,��*�����Z��w?�Z�����d4�����¤/�I��yEQ��"Њ�̳g�>n�:�Qv��?�?@��!������Vz+nB�k����ϧ� 뎼�P9���s�I���7��������@��ͦ�~e2�s��o�{�-�A�����ڴ����sX��R?p�z0ϻ����`��"q`!���Q
�R�5�LlO���SdD�/Y�
�a	`j��P�?�x�Ny������#e��w�ːB�'=� N]�tU~RYK���eZ�x����?�wPH�h���T�>�ޟ������/c�R�������<��axfd<�_�}��˵����q��յ�k��o�qyу]]ݨy��-����6 �pQa��%`^�޽�孱���&��f���t?F!�k�Me͕5!J�9���LOr������ٹs*��wS%L(�2Zb�����9p�pǀ����Q$V>Y.��
��J �'#��cUc�B��=�>3�a�ųJy���ݺ㡭6�N��3�����g�bW�G0n(�y�7Y���(�"�L�//]�9�O������~H��+
�2x�Iz~�p(l�xZV����]�.�P�����z����s���:l��t��m�1�c}Y+�*�tXŠhT�{dUQ�-���lsR����~�UH�b�T�j�\�ϧ�rʧE�L��i��[�z���x|�N��F�
���%m.ޚ�G>7�c[��[����'�! �r����>N�K�\��75nN��"�)�&�w7�����E_��<U�r����`�*A�� ����'U�X�|�@������J�T1���Bʏ;ܟ�S��HhO���<�h�J_Ei��g�� �')�/���y�駶i얹�p�s�J����!�#wj�)t7��w����m�������-P�ޙ����
��a_�l��+��<3
�y�M���O���ȅ��HH(�\tw/��XEvvvn3f��{��/Z��*ڇ�_�`�~,�;O?Myy�; ��E�v �F�:�r�7�Y��>xܸq铓�LP�tEU��˃E(�Q��m�UQ����L�|��L�cu,_�Zuڤrְq�f���yq���.��Kyq/�	J�MN����g�B�j�\/���t��m�V�*\h�p-v<z�C��l�%p銟0^�}��Ȋ<��s��3�ِE��SOn���sJ�?��/�0�̧*�W�[�gf�Y�&��-CF5̽���ho�b�ʬ� ����q �]�_�N�S+y��DQzmy?��dXN���k�O���O<����\~��ǿ��˿�ӧ�H{�meEZ�܉��s7C!�����r]^�,0�!��e�a�;6����Ea��Wm~��_Z^V�"�Ue~[]������TAO�M�>��yYm���㓲�d]���D҂?�̼(��!&`ѽ�,�^�	�wQI���O��z�(p͸�QQ�'��L)@�O�QAA�>���m�E�06�g���4ߋB�Y�lN�G�b�#c(��z����`�R�G"w�� \zO�\4�s_��%���}�q M���p����_��| �����U�<���^ߵG��Rm���rV�?��y���)h�����'�|mCC�%����9�J�]��K�4��D�ȍg��:�hk7��~�3fL�e�F�eVL������}��g-��� ��<w�)�9(gS��~7��sdZ��m9� ~�6(�Ϻs$��C�v@�����/����(%'�r�H
Yi�Fۙ�5'|ʊ�'2�zi���~P|tO�z�q+;H�,E!X�����/�} 8r�a3�%�Sͭ�S���_~W�T��p�G4��h+���kC���[�-m��ȋ�^d8�.�K+|ݏ�j��.�3k�Y}�n�<�ӯ_����_��#��ܓ�/:�gRx��!,��L&OE�宥�����=Y�\׈��e��a�6iA;��@����<����"j�,�_֢��I�ϊ?tw��y^�Τ�D{$y��M��pĔWT��]��d�+����w�G���a�1?�ݑ�v�$4�X�:V��x�_P�T�P��QO(��K�R>��9�oX�dĐ+O!�㓬��c�+ݏϋ�p��֓�c�/Y�����z��B!�G&�%=�C�א	��UUU՞�<���:
U$*�=�]�s!kY�e\娹Ҙdd�������s�(�C{j,'�A���sT4/��Mw�W �L�%��m�ng�J�gȶB����%���W]u�'N���^E	�����_?lٲe�&���P(�E�Z(�mƠ	-��|�����
�d��
���cҜp�rQv|7����wb���-mQ%����/@K��*+��s�Y�9bd,�G:;;�^�y�U�!Qc�6lذ���/ZB����,:ml�'�S�G@�^�������ŊP��6Q^����B���M�Pn4�#�5BqṸ���nZ�ƪ{�l+V�X���}�z��6TVVvvvv&����x�kkk�.qsss��7�<�����D"1�ϩ�R%N6�;ǢQXGY����E\/%�idz�?��}�dp���ʢ��mŕ	'�Tb���;]z����P�+���TC�ВiӦM?������E�L��W_}����vk8��#�b�Kg�t�����u��7+@R���h�vԑ㶩���=l e�P����Ӡi���.g�qh=C�����)P�(-��O���֯|�+����y���jmm}���	�*|r=9�f\�R:.5���)��,���<{�g]�s)և�9����Ҧ1�J�m��u��ׯ���c��3��,Y����n�<�L^TQQ1P��F@�m�P�R)))�LP����nR>�����^����I��C�6�#�S��{K���!X��V����>�Ogg��&M�����/;r��&j�̙_x��7~���|Ruuu9�� �+���L�uG&�7�u9J崓�uhS#c�y�\�6 ƺéM���V�����ZX�x�O��o��/�~�ĉ�͛�yPvwwvv� q�xpV�y�mv�����92
`� `}}��	&��\���5���/f���\�D�)���K�i��5k����WJ�QG�{b�����I�V�y���	<>eE�{��vw�()Ŷx^e7��ʮ�3%N#E�꥕����&L��ùs�Ο��H����Y�f�O�YUU%��!(�rPQ��Ke��=hs�|)v�J��pD'%���~6S���
���s�euf~�P��VvGJ�mPS�ȕ����1��a��{�wP"�x���k��/�uQ@o�fv����R�t�u�]���N8aNO���g���[n���h����d�E��Efܽ o*����\��mI5ֳ�AEe��� �:�*���������'��(9A�O*J՛H$:��˞�������:�����&��;o��§gE�E�0�:g��M 4�S���{�.gs(Sg�j�i�e���E�p�����M����8_�?���W�"�HcMM��ٳg_s��Gg��S���1���NS%(��L��<=N8�閿K��A�,׭[��c�=����|�w�q��yvuuUD��#cU��������i�lRY�/���˭�p���|�S�Ac���x�{|�ғrPFolll8p�G'k�܋/�8�>�5��;����O��������G�WS3`BWWW�F\�@�|a�I�m�P�����o.�W.�v  �O�}D�d)��H��~��UJ��Xuu����}͸q��s	��yh�%�+�1�(h+�_ ��"sn ���[���	A�$_��*풿�8��L�0�P(�p�'|����Λ7�Ɩ���*��?Q�W+N�o\HAle�Q���ԙk �2ʌ�� �έ�����O���gd�RJ!������C�wڕ�>sҨ�:�z	����n��sK�~�g�S*+*noo��!J$H��6o>��g�N����~�K�2H[�X��&+����t_��� p"[���i�a��[��kN:餜TOj\�c�<�+̯,~Q?���xBA��~o�_���;>7�@����q��{�8��C�P���:��˗W�r�-��dӧ�VTT�+�\oS
 �s��Bge	+�!��������A�G�ic�{����lR�*ڔկ،�&����k��j���5gΜ���^k�&{�=.���#V�Z������-+UQQQ#�I�-�Lv���l�&�|7�M�e�g8Qy6B��>�΂�$�������o��7��>�z���d2�`8>��� �G֒� ˾'߷'_�&��A/)�mݸq��cǎ�rG-�ǲe����_ߵ���*p��.�+��̜�H  �IDATy�C�T���>��/�V�	$v��Lr��^A�A�	��h9� ��ۦ��������:�����g!���=�͟��g���u���S�x_����D�	�BeA�Y��=����$�t56�/碌��L�l�dM�B����S>�+�r
��M&�=u�W���O��ӹظq�QMMM����k����,)
�h��+(�#�z{���9��3f�V9�1�S�zÆ�ǎ{��X�����ȧ�x<>����wSi��1�}�qf� �A�c.�WO&{-�4�S�D�o���}_�-?m�p�)2%����Æ/=dԨe�_}������%�߁�������y�o�f�ڣ=/1���r0��1������G[_���m�c������X��l-�d�+�F)���(�!zuvt�C�Y��b�!���dk�,GnL(�[�!i4e���I�?o���ow��ߞ����[��0&��x޿W��{�ҥKw(?��������YC��h�H��СC����&�Tjoo�ڰaC���2���E��]�,K�·��gw�}���9C�2g��i�������p+	�{�����[B��F��^nhhxvܸq�������˗W�����4}��}C�P�"��}�z���^YY�d!C���}��uo���߳�dS"��������(e���3{^��8����Ic�e��m7���D"������5;�Õ�}]���m��n���Vw�X���i�<�-�յ%�%�G��F�<��G���СC?�6mZS>k���R��Ʋǽ�dɒ����������6m����N$�
��D8��ɤ�,�3&	A�d�/[�掻�q�{���F��x���a��q@�1i<�Θ4.~2N���O~�߾��"a�ya/�¡d(i��ԘӲ��1&�������pg(jO$M�H���΍w�}�_�������w�jjjD�����Ӳ��pWWW����-�d�-5���ye�%�ɴ��L/0�LF��p��<����T�B!�3�L�<��o��S���z�k����9��K`�����RH3�]��u���d2�Qc�t��y�
��P�q'��L&�{�GH�1���J$�Ϝ�e4jMd��:��h[(�t����9s����px�>}jR�r�|��i��~�`���/o�{����>ӽ_����R�;]�lV�<�8�dKE}��P�}:��%�:]��ʪ_���TD������ͻ��]�0s�ѿ'.�{��k����m�lI�w��Qm���*/-��'X<��j��/�Lߗ�~N�Iw��~u����Q�G֩.�~NU�6t��Fc����q���K<"y���!��ˉ��g2ټ�OJLI[`��j���A����mP�C����X��9�?���cfAt��S�b�b��_)��%��i@k���1O=$���&,� ��~.�� PK   ���X��̋<I  }N  /   images/9a5024af-9389-4391-bb94-e3c02dff2ccb.png̼uT���.>� "HHH	�t��-]J-�((%�3)-C	*) �J3t��y����s��;�]�w�8�5�3��]�����g�&�"1!!"VV����� ��-��~�L}����;DɊya)k��_FY*�(+s��� v,p��h���^K/�]+ /H8��k�?�X)A?��;;��V�@38����K���>���LGVYxױt��vv�s��a����Ct=���,]�x^Y�����qr�[G�G�t��x������.�#���1��5����-�L��/e]ܬ�xxyx��%ܬlĴ��U�$�d���*{{{�x��ق�����y��||������|��ݙ�i��ڑ�v�t��z@\�1�_�v���db��=����#k������icJ�Oyx���6�y̷b/ >֎Fr'�<@R��"���俬i��B�sM���z��n�.N@����̿*���3���?f���R��_3)�+��� �j���3]���9� ���}�Ć'd/R�e�<���)��lqD�i���$�*�J)�~=e"�7����%��n�|ƚ�a�^�o���5�o+�I����.Y�b��^K�Cz���b��/�pu�7�
�-6޵�c(W21%��V�1^=K�w�����d��}Mc����l8������ݵ⦬��̩�җ��u�S7�/�K��~�H!��m��V9G̓ERҴ/�d�	�00d����V?ׯ0�~���)Ʊ�rs�>@U��5e#��p �_� #r<mg�#m�P�y~?%��u_�i�=�NxT��{����ƲtS�g�0�O�ڞ0�b�v����6T��T	Ӥ��%�t�z�˛.�4\��Qe��6�)�#�gqݢ%�t����`�;��:H���6`	.ᅀ��JS�쾄���>�����$<�����!���7���w�����}�<��&/usu��0�{��?]IS�9O>�_��x����c�D��O��Wg� H����A����ηZ�-vĦ��X\LZ���Ӕxt���U,�DL�WdȠZ���}�xڛ)��@�w3�Q��<@�����<��d��~�v���Ae�uu����%���XR퐔��x9�C�D�8����Hbf�}2�2 ���K|R��V�ӾJ��h��,a!���o�5~���Kq�A�7�uN3�=��
���E���sA��]��ʡ�)����*��y���+����D'���]l@'�5�y��MOL��</��^ťR��t���_��T���%F�t��ɳn��Z⹱a�Ó'�3��i/��{儹6�QI�����ɟE���/��������Ь"v
eޱ�"�[�4G6��8�i]�,�IF76z��YUS{ҟZZ���p�*�2~�1e��b�їw���wr����%K귕��U[o3�I���U0��,|��j�h3�ݔ������t<������T�س+})I����;��f����*{�T�uk��A@��b�=8X�{��j��,�p}z�0v��z>oV��p:���=|H����méq�F@0�Nl�@��riY%�x>zܛ��c����k��;�Fl){��d���o�T�K�ݙ�2x�=]�4Uk�(�� ��y���@�N��> �k �c�u2[o�P�l����2����hCP��n��Ͳ*>�|_��`�7A�j��4lK@������P�y*�$�h_+;d^����'yboT�گ�Q�G/Y�`"�١�JV�&W�H�����	�?�s�y�5:�^Y���޷Ws��(*��}s�$P�ij����?�
_`�:���p�D��R�� t'"�ra�G���]���om	u�9���j��A�nK1�4��b�wǷ�����Ԋ�m~ѡK���J�9F>,�M����w��l�i �9~q[���cQ���m�]s�{@{�֐��]`��as�`�4�����ό{^� S��#I`I�~%���3u�J�� H���)�/q�ݲ�6�B̺]¦����.���J!�q��������k�o�x�ݣ�+��iB}}�k������+���ǫˋ���?� ���^�m������8 ��������I�h�V ��Yyi�Ϊ�J�B��©7?ӟ6T����4�u�1�\~�N*���[�����!I��G��[��n��F��
�	�����p�-N�r�����ﮱf2����+��Cǝ#�:y?��	��_��U�Q�`�Y}���j�+��U�v�?�}}�P��i�MM3��?TU`M�Ը�Mb�A�l����Y`����Ѱ�J��|���gN9�1uJ��'s^b�,���di ���`j��w�@2�����˝憝r�bG��2�ux;s�D-�6}��:� %?��|������@�'�Hr�[u����i�B*��pW��K�65)un���m��]�q�MD��;|��hꆝ��,!�Ɣ/K2�/i�P7 X� �r[�%?m��K�i<
�u��9L*�b�ԾГ.�wċ)����]�v/F�����r#~�Ice9�����#�>�%<4��1
O�al�<؄�[�J�!4j C���wZ���r,J�ۯ/���A���9��^f S"��ۅ��U�g���j����?MH��S1*�} �K�d��pP<tP�jt^\!��'��\/2��qu�ʩ)� ��<߀�9Ν[��>
��d;ϲ�����3x������.1/����j] �V��4S皽�|L�����s�(Ԅ'-P�C�7��b=;�z �$lɵ�݀�g9��)��1�zUf�&�O�o�!+L�:�}̂��Eۥ���l ��D�u���&���V�BŽw�<?Hs�O����6���X�N�߶���3��-��b����{c��9�l������z|Eh
��1f��S6��髫��b��������ܼ��ct�tF,��!��͢�O�������Ő�]Lt.��R�d���8�MԚ7���̠kN��B����pAw����*y��*)80N��0U�܍D~��"g�	��>���`L���zl�pa�M���<_����_��#���/��d�|Yy_�͈uW�[ݱm�������x';�"��HjI�3���
�2�5�8��2�;�W'�����@��Hb�@������٫��)�
��A���H��ը �o\��~��H����8�/�f�Y����Av&�Y��A��B Fe��U?�_�@o�>;��s��m����:&c�����5�t���3Խ뿲ƀY�Wg�"*�
>�v�T�����M� ���`8� 
:���/6�}�����I��wR��҉�x���g �5���+�]lcit�=�QQlW`�{+�ti�tt��J(B�;x�9Y�\z�=�JC5�z��'���"s�Z�D?�Z,"İ$�V��^!9,��]�(���
l�:i�>��4��-�I�[�V!����] ��xyB���e�QjPų���ӠS�R�S#e ��H|�w��n&Z֐�t�#��m듭��v�D�~Ef�Ä���ۤ!�*y��hɈb��U������@*�Y ������`3�r�W�B4/1jhi��Kj�x��I�D�[:���q/A�N��f��&��������o
�^"RC\=ۢ;��m�Իw�C�����q��I`.�?�N�P:��$��/@S�j��Or�Rh]T���})d� ���5A�q5J�ٓ�m `M�E�jL�i�4@�@ �dA�]��?�����-p��?�����գe�ύF�T �cgVt���,�̲������^��a� xNLJ��kz3t/=MX׹T�V�6�L�Țxw�����Fe���l�M�A|_��< _
CWuttԫ
?y I�����Q����q������J��h� �כ��H�io2�Ыa�N�pa�b�G ��Dh���_e?��f���x�*��Kߛ�gzte��� d|�Y?�l,H�F@	� �℀�**w��ھG�BD����G�c��O��f��*����p��T�,A2Adjd�M!�f�@����z�^�N?n�F�k)mA�8��RX��bs��> Ow��ޫ��Wa�U���]��/?��y�����c���%1)���h��+\C��>yu~h��gk��%�n�r���T�ڛ�����ߝ�gRt;<�������rK�xd���٤hˉ��="si;����&u+�P�Ę�-}(��o3�K瑛�>꾤׵��Ƀ?��xH�ƃw8��'D�>?#��f~�qH������#�}OG���O�݂�67�DB���Vh@y����\^^�XW�# $a4��\Q�������i�"cH!��=��C�D���`45���*3v сʽB���X���ku��UR�Mk.�:��e=���|��TN��x�`E��\�S\���F�����2�����i��B[�!�~9{�>\���&��I JL%a �`����:Ao���"ԭ|ٔd��/�Ik�ɇ9�UA�H��Ad�E��f(d ��T��H��Zp�^�kA�6�>d$�JQ��#qq�TnT�w�@�Pʆ�I0qi,��s��:_I[D�)���D`�~�r*��e��goN%�c�0�8�5�������@�H]N����~/FGDCl�(�¸X�>\KQ��4�W�U+�9�ř�Y}�0Q��B��_&]�-`E EL���FӺ]�|�ٱ�^����_��,R%��g�2��ع�
� ����~5����i=���4��hVG���c�ċ�w���wf����,�+ p�������JU�x�<7G�'8�@���>3��X�6q�����G����#~��ս�ˀ��V��H�	���c��	�s�7#�`�&̲ȭ'�h$`�l�T��������7��Hp���M�ϴVkD��\�L?EN�;�A�'m�ɀݯQ���@V��������A
NsT�����C����+
m ������~JW�)�ښ)�k,�� �����V9�L�e�ص�JU5����r�z)E�{���:?��+�*8����kZ.u�Ю@�r�{�*�5/wc�
^lM�:BW癟\st�;��Mp=�5x�g�T�l��y�p��}8@
4(�{�׆�H�U����v����Q<��<� L��h�H6��Ne�����\�ɤc)�$GN��\�\��/��$9��;,!��2'l�47)��s2/('�M�{GI����*����x�+���߄iJ'2���
.�s���+������.����������(��Ķ�*�|�y]�����U:�EN{�9���VG��R�&���g�6�*	o��c����1^_��;�� ����Ăc�.f�Ga9�>_�K�N�#�JiY?y�e�U��|+2x.�>:Y����gc^X�׶,e��bK?i�����䷏�S\���|u[�3b��J;��=t×��^ 8)�g�W���0�{{�i�������T���߹��@��ǨC��ԓ2m)��[z��<��;�}x���;d"h��}u�$�i�h��7;��ѼmV����>��pv? �!�6@���R>1dLb�L���5��_ў��mVa�V�J	Q�}��ğU�F�K���QP��㴙p#��̠F|;�g>&UJЪZ�J�ۋ�h�?�@�t������]JV��Y�>��!��pL�Վfpf{����&j"5vQ���f555V $׸,H-����)��*)i�9
gȔ�ؼ΁������ht25H��$]T2�Zj.I�b
R�voh������#�����+	A9�
?F��94��CƧ�5%���Ys������ 퇵��謶����9&��1������&pk�)hj�B)RF���s��_�f�k>n��x j-�'�L��JR����y�p�ԟ�}��A��yW_����g�r����G'i�	�ު�ڟv5�cD�q�)o�M߯m�9[��t���}�/"o��hk:�������=�sU�1�{�����IG �M���x�t�6R�V��=�Y��0��A�$��}}�+{�o7t�6A:bRZ*�����礎��g�<h\&�G��b\|�����_;4�K�H?�єJ��_ʾc�&�<����{r��sKC�%�� ��\�a�f�d"ss�p0��g��ԛ[��PRu�{v�����t�"<���(?k��@n4S���y���#�����S���`�������Ljb���}m�e���4%�}�k��9虃\��"���o؂N�*)�A�H�TB��DZ��0+�)���=G�nO�ć4�c��`�
1��L��Ѿ�w�C�����O���U����}U^N�3�Ls\��$�g�C/B�;�tV5[�H�@TXum]��S�8��H�}=�K���[�Y�5ď�zf�����}����i~CE�"6�M��OyF�V���6�w"ZD�ﳵ�Ų�<��е�~<˺#�ݐm:��U�WX��a9T�+�-f��Pf�Q����Bg~+��n>�+,��d][_�
��������bO���bf�GRsu��>
��W��-O�-��h})k|*��a�\ �j�4u��������+��{�(%�n��R��ET^%�N[y�r��J ;]�֯'����v�_֍{^ ���]��y1���8�L=MK���8��p�l �߳+~��x��V�p�}k�Eԝ����{@������z��_�%���U��~��#��i��l�d��2�(�۶U?Vh!%G_C��P��\�n�ҫ2n6��ۂRmK전���\�X���Η}��V����:D	�K�)�p���W�eL�C��g(���)�%��֚��!�O�����Uiujm���u�8tl�*��x#i��2z������mr���W�#�q�Q�(�$aŚQ����N���ʽ���D�1٨� �uڽ��w�}�~M�܆�f.JHH����O
걱#�V.�с�W� �=�x��2�}��:���?���b�U����jA���q�eQ�,���Q��c�xN71�?�)k��t%��6=��>���ck��'CDC�����Y4�R5���1{��qU$�ZJjj-!���5���d��O`�`s�ҿ�?Lx?�e�<N��� Zdo(drjJ=�!�E�?"~!/O��D�O��!���ej�la����	�4�l�Vi��C��������j�6��"g�d���v�D����+2��&0{KY���	�g9Wj]��+�ug�Fpr�R�aw�^����hɡ����|!YKyB�9�_�C ؿ�R�,њ�"��ls�h�DP�MB�T?��|�r
��8�kLS�*7
U�W�+����u�rZ�cUj�������#aԫ���c}'�@m�g
�� �����%�$�+�Oa4����������^~����hy�V�@x��Wo��Nz�FSSP��0�؁2非�7���4�Ӝ�YBr&b�:��h�#~<�K���QXoT�|���jjV��-����е֣��76R+���l�w���`��� �yY�J�'�7&��sy�C�讋i7�1�B�
i�A ;b����׸��՛������3v��ë�j���}��M������V���h耶�K���)���u���g�g��xe1e׸N�5���W���L���}ɐ`j��Ho��=x\k�P�-��Z��h�Z,�B��o�z�|g�O�	&K�E��8L�Yi@��1�cMS�}�Zz��v% `huT��g}�HG�s��Z��O�/�|1�����D���g[��<ylYO	N��8��7���B��X��o&"���aW����t�6t�L�~t��xG!z��H~>U���B��"�͖\~�Մ�֧1�NCY�:/�w�9�XU��N5�E�>nU��, �x��v��a� ʞR4�|2)�Y�#�\1=�4�L~�*��y�'�Q�&��|�v0�܍\��zuҭƶ'�Jр)Wt�W�)�6^���� J����NqC�y��/�h|9<�;�	kV��}&0+��<��0�Ѩ�q�k)�*�8ӎc��.�?q�|��&�G�^�
���h�q�[�)ʜ۱2�ѽQ rЌ�𫭯��_�=<�}fR�}5a̂���R�Sޝ�5R�;P5�y��E�q)��l#>R-o%� H�N�py�����A�q�RxZ%�w[?��ii �p19ۼ� C|c����j2�j�C�3�bēDF�2�'�<$9����QXx>C�p�퉟`��$��fng6����3���Aձ��?��gڢt���a��ۺ�<��0B�Ֆ5"F/(AA`�y g����F���S�C�&�a�#�� qUn�J�9�1��Q�o����z��b���aV�E�%����A�@�i (�/� ����v�����+��W����MnN�q�n�{	^X�źM������S�SË�Jsw֡��S5�/��ԑ��ب�d�w�6��p�n�3Ũ���-|7��1�i����eQV5�g�Ř�K�n�d@�#U��x'�<�<Qc�7�1�YE����3Ї����b��6TS!c�}��W�PM�2A �@dƽ�J�hCU�GF��M2�ps��,�B �5qؿ�25V��$�oi�x4���
J{M�qȓ�����Ns��Xg-�����LE����N�!KgG�P͓_��zZ�o�vJC��07�`Eg�V���N��^.-���
�/h������8X߻vdN���>��ݛ�C��M��<6���X�tlR�y��n���'��_0	��K�5�P$�R>hk���o�C'�S�a�2��|P���MM��g�MK]=ՔEZ�7�C$ �5�����Y�׿A
�;��͘�����-�w�>CTQx�S���L�!�
��=�G5��|���K-�ް��~����[9��N�}xZZت/P"_��V��d&l��If� �Ԗ&gI[G��Υ?�Zɉ�g~��hwT����yZ��feU��f�b�Ďժ[�Ϧ6�/\G��,���;���/(e�]�|l�4�,J�m��=[�8�T� �FC/��a��PҤ��G�C����U�Ӻm+�-ń|�Ɔ��֛H��ǒ;kyg,��|c����G���L�$�kR3f�	'���Xa0�V��Y���tT��=?C5}(U&b�&��i������pv���&�p�B����B�)���'U;9L�c�;�u�i1�����$�?����^������ί88�Ki&I��M�գ�tӞDr�QǢ��d��TV�@��7!�9�w�N��3Uڒl�l
> �)A첮��*Y1��t8����K/�+vsNa>++kn��w�Vq��U���>-�t�vy����.��5��\��Y!��U��K���W1���Y������wԞ���4:���kv&o:ޡXj�d�=�´e����g��vd����������b��������������������(	r��~ֳ3�7�Kq9A�Ҝ�Tt��ig�S�s[V�t��M�s:$gה�>����n���h�ʋ���k�/p��*Զ�n�#s�Ƶ��][�:VcƓ�3��\�8#��b 4Ν`&E�u!��L�~�%x�� ���]34_u)|H��R��$7(2��(�?��̯�ٙsv=�+�g ������B\�ˉ�����b��w�w�'�oҸ����JPܦ�����|9+r�T�H{�*�A*��N�a��~�c��Wu�������Tw��z�\{u%W���{W�~�E&��cm�G��������eY���c.�p�)�K�ح��a2�nY���{HǸ�)�]����Ϻ��It~7bچ�u\{�<5�W״yo�{e�����ޱ�;(�@�vY��6�\�����;~m���S{8Y�w%�+�����ҡ�� -|FV��]�I�ѫ�h��sU�h�&�r�K��>d�����v/Bc��v��������%���w�R�m�c���~6��V��^ΜwLQ��VU���hS��!���~�Un��`���c�4s<v ��Χf�ܺ������TAEl=C���e��`Jw������g���Y\L�+m>��X?X\��'�έ����fg�o��.�_�G�h����ǣj�^,T�ΠZ]0��j�
8BW�jx@kd[ͯ�^���ţ�i���*����ō�����Ax!����҅'���_�?&3�뙈�CK�OH�N�s��.�m=��-�N�1��J.-��.�5���&7H�[����yE���=���P�La��.�
l��ڗb��_��")��峅������GKS�;��Ē�`J,R�&"�/�*vqc����Â��ieKϼ4�K���]� �o�����@{ϴd�^�i�q�Kp�X6�L4�ZR4%�D��>=Z�	Z���������R}�<������+E�̇���4�4�ݞ0sT�ˀ���Wt���:+��q��<�W�S��U1�I|�/��i��<R�2�UK��ߤn�i�:��~�RUhI��3�Z,�Z#Vd���_k�C%�5R.(.t׶���ٻv1�U��R�(��X�3��k9�=n77`�6��e��%/붒�s75���V�^�6*+<�ڄf�[w߁ڎ�Q�M\M;�Jcb�Z�=�JJY�����Z�}���N������jx ���,��~�eX�&�5�?��Z����%�>uy/�y�3y��Sp�/#�*�jf���5��#�V7-�Ț�U(k\�&��G	��-���BN{�b����&q�$s:�;�A�&>H$�ŕW��Т��|_��J_�r]&Ϲ���Г]5Μ��Wx#������Y���ע�׮�t�۹Q�S���ʱ�#��~�ɽ#ʕ�P�D�r��}F�'�DZ�7��Z	�|�8r�#��m��Qy���L�"�F�;�:�k�+�Ԩp`w��`fЈ3�{[0�
E��J;/$��8�l�(��W���B�pn�d��?A��Ϟ\�I�@o:w�t�8���@��/V~�UM��W��6&�s�-�~���}5��~Ӛغ��@L޹�Y��1~wm\We�l��B���B L?�V�*?��Cߩ�ig�N	<�%MZ�����=��}��ܼkk2��f�o���dg���;n���=YOc���G$��Re.TI*B-Β>���#�+?k��׼�6Q���X3�f����L �<�EX��OR��x�^���&h�N�/حcG5��
.�Ȼ�3�5^�۠�(��/�UZ�?�st
��d՗�?hR��9?�����*pw��X��t�vu���$uV�QuAՍ���`����\Z�V����w攼�" W�.]����ǫ��FFF5N3BS�.yo̚�V���7ssy<7G�y�_R�#���ЕմϤ@xY��*���}4 2n���V�o����R�jZ���br��v�;X x�F�9�Tx�=6Aw%b�\���; c�<wj6��^��� ������%�òrؾ�$6�p��G~ �N��͡��Ʒ�6s�,8�(�1��
�v]�'��a��	���v���9�s��%�tiG7����R}�F@I�k���=`��a����1:m�����ky�ak:�yn�����$[��%�]p��	�	n�����^�W��^=u��{n��y+]�qK�CfׄXî�k���j��Y�	S����q�`9E�|n�Jp��R�MG��ܖ�V�U<Ť+�c�"Vڤ�i�mԮ��Ƹ�5פ=l���^��'&�l���qo��:F��w��} P��-�RĚ!�y�`����_Ǹ��Qd,0�Bn��Sjf�s�ak�j�U�sL���{]��O˗Q�a�m�ÅIyI��i�!G�ݸC!�����P�h>T��{ �����&�ͩ����T�X%%�+6+j�"ɺ?UY#��v���ھ\t�R��8��=pO�0�����6 �oN�Jc@*&�<�LCOR��n����3	�q��A�2��Ĩh77*��e�w�aK[�H願6g����ˋ�]�43m�B�iZ�U�h���tbx�z����z0����ࠫ��h�=��8�:�=�_�ӿ�T�H�>x�'�mczS�"ާR�ڮ�6�Z��FJMa��� ��VN�Ć??�?�{�H��)v\�z�8�.ȟ�|��2���A~�e�*��0\���-����?a���	�'߬J �B���^�0�������r����C��(b�ߵ�b���j���,Å7�4�g6�t���1�卂qZ���Re�j՛��m
E^ �TT_�2VOm`wJe�Zb��i���|��0��z�nC\vSw$�a$���x��m�<���	��lO��Nj3�џ�$�E��I��i�!e�ZXjf�J&��`�M�`�`�0x����6ꖱ��	��p�cX��d��͏���hY#�+���^�b�}O���oD�	O~�&�c�<�)�Pz����y��:�d���|6,�՚�xk�\�	5V��|����{�qr�C���\@� 9#W/6� ��C�s���Z�~1�������
�2Z�WP<D�W+FU>��$#R�o�'X��nx�fp�V*�Qs��7P�S�,1rzS ��wV P��g��< qȆ\����AK��0`�KᅻN�.���c��d���G[a�#����x^��֞;���2���ff���b�� ����u
S���,�[�(K�tl�n����i�0\|�m�.�����)����ՙ=�*�W�n�N��/p��y��R Uú��Ӎ��4�q���A���x$'�� ��� �%�Ök��0�����N�2�d]߿��#�s���E�#�����|L'�Wѽ'�ɩ����n�עiղ��H���=��8rC��h!�{|+d���E!��< ��|z�^]�;Z-�~FL[ J";�<��]k*������1lV��mY���:ͺ������2�ʏ<OI-����>�o��A�����?�g��yafƴ��_}Iܜv��B�2H��G`��0;G���OGRq���� �����5��$�Y�O��C��I�"$df⧋=*Rq���Tx���]��������](�R4ւ�}'Ic\lѮ"�[u��_��'�fB���~���#2�����1��_�M��
�4_?W_
�ly;Ҕ�=�g-G��ތ��q�MT*��ճ <�B��v]Q�#�������{48�{"�(�r�-�ٚ^����S��D�t����L��IrbZ"�X}	��3��wL����u��+�]��]���c�-Ϻ��bg����g� ߬�}_8�QD[D��?V��'��
�x.����L0Q_��2ΦH2Ӿ��ᮼR����92������z,����8:c���ɣ,�q�*�y�c�6��e���b��\�1>ei���r�Ik�$�ר�2P�����p8X4��@�¶���+δ���M��
aım����ws�7{q�e�+雽�ԼI%\�����u*�vi��{ce�b�ޛݙS�钩>
��2��ULĥ�&���{'4���y�['i��tw��=���#���I��X���;%C���������x��K�1�p�����G�ڛE5Nߊ�t}1�}�����dyޞF�F�;�J���.��د��DT��/:=�ʈ���^PhJ����4O�%��J�� ���xO�L�<GWU��e�z�P@D#OJ�qN^2�����n�����'yL𤋮|D�ҙzߥ��ȳ��<۾I�&��_���];��Ǥ
�`�Y��S�[�9�?}���ZzD�����̮�^�oEO1>&��;bv��N}6P�������.�v��tA�_��8r�¯��ӽ��<�"#m������D��Zwkc '��s-�GO?���3�kn[6]�>7�Q˃����W٢j?����x_0��TO�"'pzT&�9`G4��ǎ0g�v}����ߍ�S���
j�V��D\�!����g3��O��FT��?R&�@�D�C�����t�KW�';ic��I�t�ʻ
.V�F쭂��h� �5�
�RU���獣"�$�+���JX"&I��_#j�h�[�n+:�;�\K�E�7!6V�4as�s�H{�	�1���`�Q5"�m ��c��L��t*d�)Վ�g�|5���㚪�#���cj�9
�Ωҹ�0iL�_�V�p+e.�Q���{�3FF A/�m@Om�^ղCI�X2]������>�ͳOT�w�NZu6ji#���Q�?�$*���-���2/ x?J��̰'����̽P2�E����&� �T2�xt��s�f���d{O��`#$���~�c��41M�wE����J��j�m|�f�6q�� �� �����%�qˉ�걋uW'�������z���2�EV�uX0B����G��tk
9���l9�`�']5�l6�,7o0V�Ǫ���6��I]iT��m�Yģ�]}�⒟@�2*C��-,\��gex���sg��h��
����Q�6`L�n����2Rwn�x5Xaݷ��) �Td�5�����0@�c���hr�۽�:)�꘽�~a�3=!�67�4��Ό���>�������Ȥ��Q���4�H�[Gu|oS�f
I�y�;��T�������!��3�VX$��`(��g��U����� ��6>B�X~��1�\�W,a���EtC�ʹ�zd�Ei���)i���S[�+I0�WYQà�{���WX������awf�)��j46?u��Ҽ�<�-�&~����1���O=Mk�ca���([p�g��E���ԏ�Z}"[#��G�FjY���OF{�ԥ��N�����4��6m�f�M_�3�\g2�T�H(��+�q��g��U�7 �ɺB��LL��./a6@�W��v�YJI�}~tO����Fd���Ѧ�\���%7P�Uj��:���р�nh�s���m��jW4���-����w�K�w昞8ZYs����˙�H��E������
��._�)�ͱ2U??�(\G1���-��n�% L����<�{j� �8����{^���4��Y�܆�@p8v��N啾f�5� ,�W�&B����U�����;(�5�𥉉����c���uJ����I�����g�W6x��"��/�C�����vO�VD���'}5�������ld��i�=l,��`����:��Ś�(�!�53�]\�S�F�C�}�R�R��ԍ%<�ۥ��p
vge*5Z��&*��@ct&6(vd��GZ̸R=:�8T�l�ؠ��3��1�����YcC����������Ҝi�(Rv��)S�iJ��rO��Ƽ��4�VH�6�z��
��d�J;�2�Թ ŗo5��	E�bk$�u�e�4���[��˷=1�&�ҿY��ę���X�ж�����*��E���eD%�b
��n�LJ��s����xar�5�(X՞+)q��j7z]��b5��_�>��������~:�:���x5�@�*�J�A�BX$���l<S8IdtP
�6(���Yq�ZF��9�ӽ��Y��[i�@�	���!-|��@��7���N�[OŪS�l�?SᏀ�)J�y�Q�J�?�0n���%n>�b��عԐ��2�Ɯ��gx����i�{+R�R�ZM@ll�������f��wj����lZ b$Y�=՛���	bU%|+��-��v�����,��/�ȿC6p�K�`p�0�LӕJ';~��\!puؘGoLc�R�8��c����w6�6k������㹑�H��Nf�Q�x��h(r�O�c��S:x0Ǚ�@P��X�ˤӜk2�>�M%����xNQR�"	6ŏ�8�L��qR�Ps�!�X�K�v-g������)i<PC�ܻ�)m&k��ޔ�����x�;i�A���yK��������Ƅ�
<�
Wn�ݥz��K�QGpW�Y��a�����M���"aa��?N�݊I�)9;;�����M�Ŝ?<�S�����{>ĮW���K_C�$|^��p�����[�	fO��>/��߾�����m�BB �[a�f�;NT�j�ڨ�����u�R,1%Eo�c��(U3��?% �7�4��`��#�ƅ
�&�3_���9C̡DTy�#�V8C�ݿ��Z�)Y���B�tBY 9�ߒ��Ӝ
T����\g�bI%��a��(�
$�V�;s��P*��`Β\!5���j���1;���O�"�[�O#����p�eM�$��Dm 1#���Q�v~�Ħɳ�OD�38����L���[��ꙓb�� 5��K��>�1���1����o��pN�s:�?�{j"�f��©W����e��Cx:PK�������~��A��`���OB!@kNx:�u�ڐ�:̹e��'F5r�&�(D��
�[ȓ홙 ^�n�~
`!�O-�&��+�O�C!S5��@�eW4���h���$�%��(�{����P1��s�=3�����@KM�B�~��	�_��;�OԿxR?����,�[��97��~R	F8@Z�M߽�{Șq�?5�{�<<{
G�wѮ����Zb<�$�=+d��v着)pi[𶞯f=ު���Ł�K�7FZ�J*�Ԫ�[?#���}:�3	�Bx�Q�y�$�b��~��E_�/�L�Ow�N�l�|Z�C�#�P/`�?P)��{�bX��:*N3�	H��}zH�Ac�I��F�Đ30	R���m�Y0�81!�
�F�.~������X���w���?�������t޿j5M��.3 �8�ҿ�
}�� ,��u����9���Y���amk�tN�|���QŹGC��qܞ��Jm�2��VS�[F�i1�:�B��B�hs	�T�D�1�N.3�A��Z�id�N$��v��`d�������������>���>����Cd�Oǚ������uT#��yԭDcYmr�Z&1��kC�z%�I�۠��A�奡:6H�	a:�`�4�����yU�΅~doJ��/О�r=hq���L�x}����V��k���0gF�%$Zܪ�L TW7�V%�ҹ�[Ăɢ�cū�d���%-� �G�-r�[�}�E�C��fW���!������MD�H������h�0Q"x{���>�����,?�*�O��J�n����{�Ӧ�Q�n�v�d�� �Hᢜ ����|�4{�c�rv�J\��a:�e��M�D��S�7o9 ��z�(���	��%��tl��ü������d	���}��/� HВ�t����l'3~j�x��k!T����t�&�޺��6���x{!��)Y������]�K͋r�������6?!b�1}�y��\�����H�Y�q�TA����g�
G2e�J�ܞ�lmN��|QD`�MQ��>ω�ќ2���jX���f����%�9v���y�?��]��.T�$5�+��r�[|;"�k���ό_��&xC��!-C����I^�{5_~���\��+�d#|e.��t\����>竔�A�[�}��i�����s�AZ�И�27���b;���������Jcb���et|�>�mЃ�^��Cފ+��-,+�݂����JK���.e#%�*Bw�O�
��6�k»(8��ѩ@mB�1I�	��a"�Tv|���zT��0�?��=���|b��D����~���w�C��nɮ �AT��ۋM���U	Hb;�m�X-�̀���;��y����Gf�8۵MU�7�s)�/��t�3�N1	�뫛ǕZ�Ա'�4�:�d��ߣ����6H4X�+�
���d1�,3UY���dh��B|����<n�o��2k�`x��IĻY1�	q���C/ׇ�]=��dk�*-��[cf�F�#?�y�F��Y�K�>�	CYq+ie^9�<KV~�[�{ol(0��_��e���PZ��#g-~$��g���y�� i�,����g�u����t�(����x������u�(X��-�R��j��f-�y`k���Y:M��W��w������Ǩ)�;r������ʳt�����'��P^d�
�z����h�]0�#_Þ�d��� N�aW����J���!�5���/��i��8��V%��LM�4TD�mƓKRD��6|^��'�6�ف���w��6��n�y�����p�'C��g�jg��P���tBx� #lB�Fp5���aEH�,3[�(�7�h��j��x��g4b˗y� ΢ݗ��GAH�	�N��Bk�'[�/��&y�T
<J�7	}�L��;;�Yxi�6+�VDg|?
�B�OJ���O���\�ܦ��t��&+��;�u��~7�PK   ���X	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   ���X*�x}�/ �S /   images/abeae39b-2976-4cf9-8094-7a1fdb96bbc2.png<�u\����&�K	i�etw��tI�Fw�A$�4����
HǨQ������������w����y���7�
x�)?x� OIQV��L��Xi@����L"��j)H?(��z����;/��}����ùI]�+���E��K�',c)h/A��Lc���=L�J>�bJ>�'�>���Lr1�����Ϊ�8Ƅ���Z��o�3�~�H�;8�'F�"��֨0�H������+��������g����_��(kbN��q�ww�]]X���ۯ���F���K����w����;(��id���,__������E�����ꯥ��g�ʑE,�br�rUe��p���e��m������6 �J��Iec�6qR+�P��War4J��ib:�#�JhDY�ɑ�_���_�E���q�4Y���d??A_��? 1�,���0����S�8�U��VS�_�+�d��?Z8���yħ''o�&[i7��k֦���������aaabY���7sSSϢcb��ē�/����8''n�P@��W����4�R��JA:�#��b|��Y�٣yt��Q�����I�ݓN\&;�L������c���������X�X:v�"�wXn����%#A<��e��GDdh_`O�E{2&}9�[��<c�"�Ѵg�=�o/V����Iw_߮{���:�0�d[�m��J}��?��EBE3�y\é��3tp����Ȕ�̈�U/77�aQ" �v\#���Og����6Q�<�jĀN ���p�i�#�/� ˌ]��}�%��Y�{=���*�Kkb�}[�*@�L�����0���BL����K�_���Pmf~�����uG�2��$W�|ɓƹ.
,�w�Ï�%�[m�?�s�^kR��5?݃FϚ������h4��UN\�{r��X�b["l�r�ZJ�Y55��+=�|����Q� ��Wy|,�ZvH��@$�b���DJ�ca���4�8s!HRux���ً���RD,'�+���
<;������K�J�Q	:�(ǽƑu����9�j�����7�3�sy��x3�PZU���j��7��~l2)�<h��X�]������׃]m���d����c���p_݉\�e�k�nE�W�����AvO���q��~�{k�:?T���Q��Y�ߜ��W�^䢟�ȯ{�S��4D�'nk��@&��>z!���/�ȋ����´e���e|��T������$9暨�vԂ����XA��;0��TD���z�U�RQ�C ��M	����0���4 ��|X���L���C�+��F�W��c�M�Y��l�:�,�삸���+�|_"�GGG�n� ab�8B98ֵ�/���l��K^�kW���^�1��t��B�?n� �����`�·������r������g�x-��_'+�!ސHN���QbX���IDc��c�P�uj���(�?��^����>����2��Y_@,y�����8�3�WE�(Q�s5����>J.��.Z�{�u����G��Py�Z:,��:6U��ؐrr���r~��+�8���W3��z5Fb�ѓzq<&;}v�cT�!��zߐ��_��ģmq�,�/9��@2WV������Sx�Wŷ�">��_6�Ψ�ǫ�̤Q��Һv�GR�qƈ�|�㿬��Y`Pi�<?=y`�oOECcF��/$$GB��^��������ml>0wA,��_g4w�Q ���$��7訸��/�7�A�W��FT�i7N�i)*�V�Cҫ����@�Mf೟��b1�8Zu-��QȤ���������_'��GW|-��ú`hˇ��uUR��鈖�_�qM"M�& �z�
KD�E�6t015V��ҚVS4W�2� w������+}(��7�ü>���T�1�Z���Iۥ@{aX#}��������4oPg=���4a��?#�����(��k{l���,F��ܩKv��=q1���v�wj�,�����,L7e����Y�� ��!���a�n`���Z��B�B��OA���Ie��3���B������;/��J�o5l eO��x4-\{r�))���_*暹Xej�y-���TQ]�[o������ºJ-B�I��<N�,�R&Ed�Ӧw��Q�B���V��f��3�q>j�9���Z�G�.]@�#�� �Q��nyYyy���D����4���]���H]�tEr����4�?j��j��G9 -Wj�-��W��<�����F#i��`��`�ZB�?S$\�J��}f1�2�͌�XJ�_*b'��G�f7�'V�V�L���Pms�;�����Vb��-�&*��ɱ	�U��*S����"�wmh�U͂<9F��2��P��e����0�0�,B�	w6t��Vm���D��M#�:9&<��Y�	s���\:F��8eP����v��HC��W�{����QӰڃ�>*:=��ۖ�ಳuJ�7B��z�����1�+惯>�C�����Jǲ&����rB�:�=��H��M���tyM��t��]��~d�w��;�~%LR[;���驜�%L�$�At�7L	�P#e���*( ^U�Dm-QFİ/��(��K R�2�m�htخݏ�̏��#���X��ɧ�̠�@ޢ��T���F7rغim�j�y�=�}���sz��ޕ�p�ݎ\�?6�g�UJ{�^ㇼ�S�Q}�g��Pc�$�[fK�2�J�x��N�|���̞J�.\�����[�z�}����~E��*��Y�xr4�2�y^�)�&���=i?+�s�<�k�X��#.i�)E��R<�ǫo������C���p靖�Z0=���a��$�-Iɓ<����ޅ��6~���ȼ)W�P�b��ܟ8i��q1������������'�q�kkV>-�\Ymٿ~�����xՂ�ME�y��F?ž��-K[T��{�L;����f��]���OE��� P�D�v�|-Ŷ�+�(Of��w&�0�iK������Tʕ�`lK�t�n�ǎ"��G��Yޢ�K��\����>���p�,V2BF���+ʶW3����qt�]���Tn����s~-l9�FTG�I�[ל��I�ld0y05�����T}1�hy`�=Oʶv9K����ñ�>�"4r���w���[��o6��ub.4�˕����q"�,��y��&�V���%�{���w�����Q��_�'6��I�5��e�:,%�ޔʟ�<��mMTk�Q����ҊL�`��҄ti�dڠ���&ׁ�q�t��3�/�q���,�P�?XJT�9e0���x���=����߯�	�.�d0�Am�g_�{ԾU��r�I��]9!7�~jjh���#�Y����$}����+w��/_�D��G��ƕ\�6O��ʉ(��<G�gX؃�
�,���w{�!����y�Bi��֚� $��E/�SQ=VZ�0Ryd�p|!jHo|�
�����B�a#D��ye������8I�����m^��X��?9y��>�*���".��:���ȦuFbT݆��?$��M��-����40��-�4ԍ�	/.�tSneؿn:�Q��^�ar�'	J�X���M��>������7C�B��fE�󲇢�"[�c�3��A������H�2�-&nTɐ�8_�A�/��c�G�+�G�KK!���.�\��3'���CՎ3�`��"ݩ�jj�β�/�ѩ܈[Yգv��BL���x��"27�Y#�VG	�rr1 �?̱Z��c�F&�t߆l-u��m=� �:�׎h�ѻ��9D��c*� ���4�T���5�	g��8#	�f٪veJc���p��}��%���Ր��ڳ��rjK8� H���b�E'@��ؕ3wF�v��QB��d>�kW�b�o�p]�f���	vX��1ŵ��܀O�%gč�O�L_�E2Z����mJ�U)}�Xt�?V:��
��p�/�%�w, %���w�yO���G{C��������e���F�:sK�Xob*r(\;5����P�?g��Eҭ���}}5��Ͼa�~�JdP]���h^t�u�2N��J3 �4�1 K+fs�"k%ֲ^�d�����+��A&ȟE¶}Z�|qA���f��	�O�a��+���!B�n]:����`�E�?~��m��Th�u�y}	\i]e��|�>��߲e�*���[�fZ�s-us��-�_�l�?�����հ����2Y�6�U���{(�p� ��.�s�C���)�h���O���j@�{��!�^���.7��LS���Ox��y�ݭ`�����v�4��|�k�.�$J�׏���gωx������H�}=�l�R�!�fr�L�	�dV�"�6��F�NN'����[[5�'#��G�|q
��9G��Tۡ�YH
�5��!?Vwb���tx���?%A�׹7���	o����k	2O�Y*Q�р�`���,!X}щ\�d=2�}�rsf�i�.�p��p�Gq�(�/v0S�;=yǸ���W��WZD0�￲|�`�t�p�c{�_��G����J.C]nڏ�[o�f\��'�Az�� ��O�x�Oi�۹%r�*���o�\��*��e�)lV� ������K�6�5�vn��� �`"���V��Xl���'~��Z��9|���� |�i�0����0F��?�h�}�ޯ+�hM�lb���hW��"X���B�!�{�l|�2�R�r��6[Y�D.���Ƿ{�f ��[Z��Z)�ù	%��V��-b�Z�S����NM�(��nkCib���9,c8�=8Ĭ��Դp��m�*��pz"�k�����A	�����k���q�R��5-���l?mg��P��npG�����x:��Ȫ�ë?���|�aa�����0���*�󝟗W���R�XM����v�Ibv�7�j���ݓ���>%��A�f���XZ^�&�5����GQ���@�l��'����r3ՙ=�Xg���s��ʩXW��|�X���X����=w�����̻��S�q  
>M����+!�M���p�M-�~��Bil��@n}�>q�����	a�6;�X��?$�T�?t����-��[)�?�vv�Z����;f\n���g�F
Ѹ��n���B?�ydeI($s�-��o�P*�`�e��W:��<C��b2�鄧~>�O����)�B�>+Q��A����L8Zr�����,n(��|$��*���E�&��U�������?��]��HS��wK/��M��G|��	'����d��2$hbG��hot$��d�}1僬�l�\#xl��*M�uH�l�
���+����+�<�np�-��%���қ�HX�M/+�ߗf>�81|�}�;ӑ%�+V١���@����NDY=��'��3����r�Fj܇q��*]�2=%���d���]��)H=SX�;��0���#>$�W-�
=�y�{�𫻜�B�n��L��~H��T�	���^r�cO�Z	�v;�3��X|=�������K��"��� $<���e2$�m[%��P]&E�pkp���T7�"�>U�	��%��ʹL�H�--Ѵ�_�LI)��Ֆ�������#΂�k̡͹�{��Ȳ��Clj1��а٤c��-o(���ߝѺ����
#�a��qȎϟ�.>3���;&��ہ�&U�����#Lx,.���!^,nu46;*�ӝ��$*([���9s��v�[_�����9P�����F(�e2k4�h�}��¡܋�S:� .??֊T#v�zLB2��j�"5E��"�T`�lk{�����.Ҋ"��(SCx^k�:�.�Q~�7�ycf�BM��Sґ/����Ґ��@�2U�j��R�	�I9I�	k��l�Oi��� �Z�?Y���
����s��YZ�g#Y<� fq{V,�.>Y�O�򥓂B�UU�}�@�Z���Je�}�>@�/~�*�su�	��NMz�3�,aWk!�E��P��c+���)�1)�
��-f���a��k��w��U	�%�\	i3���r���:���쯩K8D*$�zy�1)�E�l�\��N�#�K;$��{ml:��ůR������5�/�ӭٱ;��t��4�I�qLKmپn��f��%W]�P1B/-�Z��e�����������Y��jt�ۿ[��J��^�l8*��1{��%��.NmϤHv¶��I�n���R
����k5Z�m�z��$�òв���r,�Vx��t�6di�K��}���ᘟ%�h�M#��K��B�{F��W�=���"\q��\�jz�NH�K|�n(��s<��dY�(�&\")t��"�M�g~��w ��羞��U]������;6���2���{N�]��/�&����  ��Q����q�sd�V�3�^�8Xs�p�:JN��t�� (7$	/��qj"��5����
	{�����
��"�=�O�����_N�m���S��{�P�T�*G�����Zf����7�e7�#�q�َ{�j���e���z��� Dڀч���B-RpE[�v����m�IFY�6���,�V�C�Lqwa�_�1�#�x�?��b��.E����ETyY�qx���v�L�g� �k��{��LJ>Suo[Um@J�1����˕�g`~��٨�oUX�;���i�)���!� �s^4���Oz�v2֐���32��ٟ{s?~"2{˫�3��r�"v����bB�|^{0��,�_$U��FJ�U����kGGd��ѻ��k_~xw��k5��xN_Ɩ%�g[,z�s���g�Eֽ��N��)��&r3�-�3=&�<����������]L�COA������]�Mʹ�g�O꯰m�/��y^r��̐O���aF	�j���]�@^�O�hj�*���2�/�:/����U��l@�9o����.O�i���Z\$��	��-����)�T��	y��[��E�}��G���Wf��pM�I^�_��KF�Ҧ��[�%o]���Վ�"oU�����2}��4p�k-�I����44�WO �l���V�؋-�z|(^[r3�z��q�ntP�0�ԎL�@�}�����֛'�5n�Gd��3����3������Mqm��v�6�߭���AI�ie��r�������Xُ�������d�DL��������<3��2���a��񊟑i8R+�1����ˉ�dl�UNHt���}�;���MӸ�+z�hs�h���#��>�5fs綟˘�f�&9`o�~�^�ເ+	�B/�F�3_zd����"#R��Dn�����:��,�ǻ���Fb�r4N =ގ���HN��t72�����5S���S��[�-��^h�x��`�9����z�=��V�����H��-L��,YwG�\[�����;��w�~����jX��4�E����Ҵd��R%�mn�U�?�B��a��@��~��b�P�#}�[�|M�}��}�s��ԑ֯_���#5t��"'i��}�����������ڿ��N�|}=�"-	�����*��VQ�Z1U�K���
�{^H}�´�xcx��m!��CRǁL���BV�M����߄]�r}k�o���@��':vC�������d��y_'U2Vv{WX&�M_�"��:�	����|���}��A��v�7�u�X�ٛ�j�O�:p&�u+I�.��c��M�u�飨f%�M��.��9C��'�<�]8�9�kX9��v��=�2%��יԁ\��N`x�3[�#�����8��7��֍&�TT��3R���ng?`:�;�f������(��q%a�3��!�����r��Sđ�ʬ�1�`t�}Tl6"�m"1{IR����EΡ��.h$|T���6�:�-3��������v�;��j����&�t�V5!��ȨUA~R��˥�b�hK���h��bx'f߫C�Ҍ�-Af�#�FG�¬�`Ix�lV�&R� i��xr�;�J_&�D�M\��� �|�?o�o-�+8Xd�*k���B��S6��S>��� �cHs��HN����^�'��
ٝ�{6��E���+k������%��Ecso���=k:Zfh������'���N����^�$���|�;���|���/�wʊ���u(�y��!��"�-蝑��yp�u�/	��AG��S3dr`��EV��ӒOAJ;�_5h��9p��	h��lԨ�t�������������?T�g̭p�J�`� ��6�/^�.�S�V����)������.�
���;�ˊٔd�����u�8��===�!<����a�ȆX��ylи���e�inJ�\���w	�R�g(򲲊�����;h#t���5|o�I�^|r]\�=a|�D7�ǵ8a~O��#(X~��5�	�ؒJu��(Iˡ�N�&#.�3+��&3��4��~}�g?�5fa�oN״5��@�;���$�>]�GX�,{y2ԶoI��`z��m�T��x�H�z%e�%_����ńg%G�}�e�����H��-�ӸQ�)��2��QP�K?=Ԁ�)�©�Xx����L�w]>��̰W1�ď.#\���W ���'z��>U��/�����q��3p�qڹ�a��^o�P/��˹�	�2��-O0INo_T��	�X@�r��1�s��T�A��G�G�H����U��t���1���Q���Y:���������(\&<K�;�.0��&m����" L_�������lt�P���K�ő�ڜ������� H2�q������써B@��<�Nv��@Hl�aǓJȢ��ewfڢb�ܦq�Jf��N"<���1Y���Xڱ�I� ��"kl-�UQ[�S�h�@<IPΡ���w_�E��"�@���R�}��9l~TO�ĴH��b( ��$"�s�\L���y'���y��%�"��%_P���c�~�8�؎S^pU)��埝?�@�/&�&{}��߻{�TxA��7kD>�J
�>�,����xGpJG-�����>�M�L�J���l�➏2E�� 7@N:��7^�~�=7Ub'�<���С���܂�"ej��q5�!Yb�]Jj��F�5�}�>!����6�����F�\�&��r�~�ņ�B�pj��M%�jT�,RXm�s��x���a����_M-+)�}�FE|�%ڞ�koZ��⎐�#U�!�׮޽��5�<b(-��p`~<B��@ǀX�)��z�(X�z��lO�����Tw蟄ވ;'��1��	�ްh����@Ӯ^A���t�ՐL�Y�r���9+nd,e��M�����m��;!� )��
����93-�d8wZ���<�$�/kH$�kbr�������_�|!��XL��d�7�	Ap�QH+��]&i��HzN�}�}=��ER�YXq��ݎ���*��<k���	
����ZB)��l��٬���g�E��	����2+�] >!�܋W����?51x��`������� е49��([g~=����~�//o�Up	�̟�/+rΉ��Nlj�m�	��rR }a�ؒ��v�S=RC��POM+�Wt�\��O����8�;���������sGG�(ac��h��N�� a����7�,V�|��&�( ��;���F�ռc���ËYV�����[� ���oX���ytr���zy2:n����9��	kĜ�F��I��El���
��� 5��N��6�$'ba�k�� S��k_�&�@@�\B�p8#�M���[�����:�9�7������oE��h���.@��2e�:U��2'�?g����4����Q����֯�4/K�D� 4q��N剌%�����pB9(��L$>]i��LPV1-�)�'1]|/l�ι�{ԭ�pGox]�Ħ��.�F�sD�w��G�F޺�w��y�~�� ��=?P���"$�q��@W�\	ߚ�G�+3B�B�z�`�����R#z�����f�=drr��u�;΄-��v��9㴔�����D�&�h>��=<S�Ш���au���6TEatt~�2[ӾH�k�u�̆�z�h$~�:L��K�L�	��֮-������ZFة��끘ʽ-x����m���r�]����v@�f�N[���=U9��N/��=�5e��o�S�R�|��$�y4�){���H"�|�o�nX�LA���[ʌV{W\LeIE�F�Ag�B������¯5K9��u=���޾uC��1[떛�Z��t��80��s��-��Qn��x������p�]�]+Iv�mrX(0�w�'��heX�������S���ș����J�ím-�Tӫ����ikog����O��u�9>���<B%��<�����J����Ux�G2�玎렶�z	�d�����5Wՙ���7���p\OY����?%�9l��J,,&)�V�7�h�c?�j���V@I"�I�$-���C��������ǁ��L��d ���?�Ģ��&p�]�)Ԩ!�w�K��g��?<���\����p�l�$o���<���=����x������f��z�PCߵ����Cr�/��T؛�s^�(�a����h<��s3X���wT6��|��&;�\���mRs]c�Q4-e�2K�p�g�I�[�^Z�����h�Z�����Z��\�0��$�v����sL��ۂLYf���r�?�ST��v�
If��ܦ)#;	��\���ӓwo�x���9��L��Ri�UU�W�
�#��-ݽ���NH�ʆL4Zp���-��R���	���׹�
�I�}<01��st�������o=m�����a6~�w��;h6d�y/2�����ĭY�����!HзQ����2 n&x�rȕ�dX�����7���VC��^�����U�q�	�˕fkd�Oш��<07��
��5�5���%b=�7W�d���;���zm�z�Bz��4��H#�:��|d#eh�sTq�ظ�?�ܸI�)']�JHP���f�	�gv�W��f���`�mXC�"X�K�Y��R�}?��8�Mٝ8����
�IE�Y8e��Ʈq���nM��:Q����mp(e�/��b:�~�D�gJ�^�;��NT��7�m���s�D�����L~��u�N�v�(,����� �;@|�~���β����$a�ɟ\"��V�5�"�*�Q��[v�X�q0[�n�GVzz��݊jә�q��� ��J�w��?r�gs�J�
�꩷�h�JF6*!�����F�s�t>��y!e��ICm�Ƕ~`c]|른�<��<��O@�C��n���R�ܵ�uH�DPg�&��uv�� V����F��x>���>�x �2.��U�ؠP��BJ�8)~ �\p;"?�Tс�g���j����4^�����!��ӝɭ��¨�\���2�W�W�����a}��u^��`��^\���ݧ:�~�\�����HtEk���e�+���P�-�������� _lgEv�� ��g]��l2oAVt&� �����!�5���E��?H>��Y�(&h=�H"u|NMX�	�'����,�&�N�w�U�B}"W����32�g3�,^��A�F��(.LR�ݠZ>D��Z�U��jp�m����_@�O�p֍{3�GF���\����dd~ĝ���A��&����d�7�8v=P4�)� ��j�in���B��u�ƹ� R׉{m
M�M����=��D��?n�����R�w��<
�@W�7��̆�g�c^�x�ĳ���;Z��CZ�(B��m�{�^�K��8�'��a�,?��XM<l�|JƼEgu B2&���#`���H`��}m�\���By�Ѓ��d�����G���Z���V}[QB�����Ѱ0��y<哈!�EVqPI��<��
����}ɟAgM�Ce�4?���_��k8�$�V~����d�Ѐ���Ce)�=x�7d�Ō����C-�@I�q���B� A��hk�.�̸C��9����8L{�e�Qu@V�j�|��3�
�>1�)6?�nC
�X�e޿�M����� �S���g��7��Ƃ�%�J�r�ͷ����M�Vd�ћ�7�W����Y"�SQu�u���B߲@|�������=�x8�
a�ߒ�aű�r��{!�LJ:���vV�0om���r>�v{���;�v�/��FqAb����  �ؗ3>7����c������Jo!�ƺ����rC�@9}f��y賗�-2c�s;�
����_By'�r�¶�=# /@�-sAt�Ԙ�m��L��"E0��d���ր|E�6
�$�U/��݅���MP{}}%��o���)����|k��6���ԍ(^l�S��w� e�����O�5��O)��%�pU�Ng�x�#�]D�e?��[�$No5ãT%ϡ_!���I��O�Ռ5a�����c��G(�v���J�f�֎k���T�8и�w�^}��#����^�W�p�uspٲ���_�R�?����F��'c�0�#ˆR.�1������=����"Ǯ00�����V�c�C���"z�����x���Cc����SL�ߊaq�g#��ൈ��ޠ��������Q�j�%m�k��g���m\C��a�A�ݑ�H��T��B�ryq�c�[�˴��#���[ԗZS���2�p�s��C�x/SlϷ������T�5�3q���9;ǿ-��'֞� �olrM�ԫc��%J��)%��@9���D����̱�0��7>l�|�fZŖ�x=��m��s�)��z�W����|Lm�R�w���{%i���꤆�f��l�nX�������2N��=7��C����x���1HU�+�k��!LjFx"���0�t{�I��/!�6~Y��)E�}Z�6Tc ��;<���]6}�1,$:A FU&�O��B?2C������A`��38����tͨ+�^1�"���qdjꙚ��h$	��?zr�i���@^^>�q|��A��E�W�H@Ys��Љ�˄ֻ+�3��-� ��V����\^f�t�����ɇ�JŨ(ss~J1;>#	�:)�(j+��Eɫjm����)�qϟ`�7LO�ʒz���ys��d�R~�v��	�\�X�	��p���7f���0&
>�cQ��#��J�a�m��Fe�\���,��J^F��2�b��Lj^0Hm�1�0��I~�K/|sv�oX���P=DD�kqܽ�p���M�vw�-,�(sĨH�7��e.��7��.�Y;��C����/;]��Y��\:%ξ	�z��j]���0����.�L���P�Mg���m�o3`	`�G����s�ia�9h��¯����1�i����n�z�2���"QAu/4�w%^ѱ?!����nS�=4K��-��EV/�i�/�@U{E�u�=������Զ;
����a�>�\�4������̡,�~��_�ž8�Dق�w$WWC�W�OM�\��O���7!�����=#��o�1^?�����|\�
���l���1��$�d0�:����r���U�e{�D{�IYw}��_ȮLO���N���4v�O����[��j��>.��e��Y �����sި>)"�EbhKK�ġImu{sNE}�ٙ��/(8�.ae���e

 ����[��"�)�=lO�=��o�˘5��?���~(��o[d?�� ~� (�����]iV�)�(o�A�ٕl�*��Ax3�ا$}�^�w�N��>������+�b��{��=@� -o�󄠰_[� �⃹����g���p�TI�<0Lq��\)���8i��{M���a�iabf�����*m�A�q��f��~F~{[��y#z{�M[�5����˸T�$���HrY��u�vp�_�w�rC��}����L���]�G\��E$�5��|�
+ί�r`�>�p�>���kڭj�g=��Y��χ�Y��<_�JS��״����'�ŧe�Něszq��}��H� �����O����{R]�'��Kp�����hƊ��P����s�I�̆T��f�x�b3��D�:���� �a��(����(f�HWWז�m���m�q������<�Qأ?O=���L���!��d={�+q�s;�"��UW�zP�N��⛌;�4��H*��YJʍa;��� �bG�2��K����>��L��|�"��h��QT��,�]/�u�^0d[hW�Z�Ŏ|��6����}{KD��Ϊڊ�^�rI�`������d0Uzi��0������I�6G{�j�t��fg��z�� ���t�щ]�~�V�Wn�n�*��( �Q�/��E�����mW��P	��2> Է��yS��	��°9g���1�W
Q�3Iۑ������t�oFR�'.���?䥲Ȍ�o�Gx1�;1�9���{�XG��Q|��ŉ��슩#X��x���KoA�!���/ҧ�� f�u����Z׉��6�u�Z�#��܌M�{C�*8/\ac�G���m���=4n���k��|��������*@�@�L.�_�i�e��O+���v�I�R�r���dLRoTp:�����O0���:�����<��TɃ����\.I	Rk�0�0HsʩpU���M�����:�B��I��FcN��q�"�7ߺ�c����M�#�@j�Un��8y��<��G�Q 2���1a���nã��|D��VJL�/����׉������Y�7Gd��hh��lm����а���]��El�N��F���'�A�xx�(r�<�W�	q�%I���sB�zU��4HD�p�N�虥[�|	 o���7�+ �d�┡ҖftpM��a���C����P*��(KLg�x���(�u]��lp.��N�|M��Fu�	7D%���:��+�I� �t���(�w�BPr~C"���)���N��Ij��6�c)�4��� Z��_az|��=�"9�n�!X���vNd���v��};~���v4y ���V�� ��F��ە�\.ǹ�X��m-�|��;7�D^O���hj�<�7�T�|XeR�8i����!Lx�j�^�ȣ���[���-9�>lis���Z�KjާݮT�����}B���Y.~{�����S�4S���	����>@��n�}s�6_��J��]xDI��x8�w&chhX8X�6&C+��X9�y���b�s���F�V�!�.ՔO�X�+�?< Yn���hd!7�P��C�?a�KV�HN�{+Woa�.:�3򞫰13�I��$|���?~���P���������b� $A��>W���92}����5�w���s��Ox�e8��d�,%�)�-�iB��SRS-��j}��]�g���lz$0�L�e
��	�w�d[=�=���f�v��������[6�
d/o�@b���c������)�f��W?;�O�X�H�mI� %�l��߱*���$����{�F[<���h(eĜ2*P�IOd�o�<��>�/�7���ܛ%�*�?��(!�WԜ��m]�9��ā�x�e��	y�T��&\l^�'1[����H0!P��?�q�=�"�#8c`k��
� ��{#��������	�����Np��`���TN�"IJGc����^P�V�@{ m��?@����.������9OzF�g �����c٢�R����Z�A�HJ%j=�ro��[�0��(��2Ju��_�z���я{9J_�������.c"��d�|��/�w���F���m�~�Lg)h�A�=\���N��	��?3�4Fg?�9x�����������i�IMO��F�c�ϟ+�Ơ���6롬����ȳ��W�VУ��Z��=��'���i��������z_R��Fu�<��z�����~:0PxY�*tV�|8����G��NT�/`�ߞ���S@C;�R�C��i��������gܑ���:�a�Ԫ��˄�k�eR6YZ�KHl����i'������(��?��!tŵ�졠�V�#�a}��P�F��ʤ����sa�I"%;Hy���vN�?�(��\�>����(������}j�v������tCd!'*�s$~��HނDZG�'����Q���ӭ��k�ç�n��"���S#�v���f���m��"�l���nO����SvC�o�e���/�y>�{ls(�J�2��gT�
I(��íS�,��*$`�bQ|����D&%�-7�O�I�Q��mE��f��{/i�<���3�QO<�W��?��L��m5Ե�B��E�D3��%���vl�M��Ps���}����а�����&tM��yؗ�wi4��6
���5��\Ȝ���'P���ꒋ���z븨�'l�WX�FQ�K@A��X�� %E�%D@JJ���CbAXI�%%��Zd)���Y����y���=�̙k�k��|�(���ԇ���8��0+ix\��i��9���?��f��w�t�^�����8�刺5�hVJx�}�Eǳ�7n��!�sVjR>a����'���ύ�H: >~/6H���4=(8����+LO��:ٴ�(���Ń�+�_�@BB��M2��vz�m�
G���	7P�zz���4&�b�Kf�	�J�ꖔ�!������"��ф����L��"j�����Ui�*��C[���L������WI�Y���[����u��}�c�����4l��3e2)Bn��o�����e�AA�U�t��bd�����z���'.����O5���N�rv�X,��ٓ�E}�ѷg�8��DF��\�D]�O|����k���N\�Z�H�=�8I������(�!�[���L�WVJ
$�cP�,�~8䳮��$��'�ш�dN�L�BJP�IX��9%yB�԰8���=`���]�~l\/�D��~����ڿ����-Ւ�WLM�O��)�X���˜|�C4`kN����
O��,H�� f M*+�����>�d�`0�ey�L�8��/��IJm~~~�Y;��˽ը~݇uW���:!�w����$�`�0W�z��lb�OOB��Z�2�y�Ry�P���ϟ�)�} ��Aŋ3�V uJ�A-Kj��t�q��W���`F���Lmi��C��]i2�J㯝Cd<l�`��;(4���K]�>/`%b��pez@���?ڿ(��g�E�ؘY�Ŕ Vy�Y��ҷ�z�`�K���w&��җ�H2ꮍ�aS.Hxlx8�ezʠ�5����R�����Si?�O��TM$Q�B�:
K�R��`V#ze�ɉy*c����,	�PH�o�W��ѕJ�@��%�`bx2k�}v	Iq��ד��U�~�g4=Nq�?�oS��E;P�Z'��(�}s�����ϗO��1�ߴ���x2e���+n��;J�;���k�b(�SK��J�%{3�v�Qv\���VI�$�#��6��J+�Q�y��١���(?��`?�Gf�T秷�z�	;{��@]�?6D�dx}�B,�,OW���.�cq?���|�� v�A3i1��4*�/;{�Y�ON�v�g�/�?���EA͓d�e�tW�ؾ��~slH��o�a����r�"�m�X��?�a�� M���'=5ϋ�uU��l�}�]���ۋ/��hk�4�	G�U�w<%��#�l�������vo���IMɳ��o��w���fղۍW�&�o�#���u��l�W��e�'k]��2W3y�DqH��/���M˵����Hƕ������}�AD-�	�DD�
�C�X�����-J��6���
�7�<~�o^��3q�]�p�%�>�2�S���'XH�MH{ؑA0��BJ�z����ڿ����:(!��8�>p�0�vS52�`~�S5���Xvv�
)x���P
)tt��Sq\��9��7k=�8M��#$�8�(ֿ�~J�XM�#7�*�Β���L�` �α7?�ډ����ͳa�a�z�Z��} /W��Mg�f��[H��f��<�Z`�j�V�䖈T�T�V�qE@�R7(���x4=T��9T#���\:T��[�^�suo�]~3��L'-���E��)�2��w�yMƏ��koVeܛm)S��I�6����2��徵�?��4�᳸vժ��m�0��I̊s}q3�8t�F�g^aOL�B�½�g]�>��m���HӢ5kq���n �w3��	
�}�0?"Z(t�`��`�f�BMMIa,�G�����x-�y.-�8�W�S������Kn+ ���7~,>/���!��x�Ә�u�5�%s״�����i#��M�whA4��X�;��!_�"�? J���G��)�TY!/�5y5_�,�W�+�����_<�t�+`�X���9}%r�R���S\�Z�]若ǵ�
��ne1L��닸�X�g���B(�+d�Z2$TZ�ؤK����9�:�h��3i^��z~TrW�����w
�>�����TcOtUgT��G�����	��=�����_}�et�ݧ�ur2��4Xa���e��b������<�=�x��G^�{5./��ϫ �`��\a�St4�	rA{�#���
�K��C�H��8g����.�����Jt&r�~w�]f�ާ!���h�9dŠz��B@d�[Tq,�)�9Ÿ��bG��`�M��4*L3�G��v�y�ĝ�lUq����^�c"���mQ��`w
2���:;��Y����\s]?Hu{�~�'�ĬQ+O�sAO�[R��}m�y�$���i��dM�4�T�g9���m�#@�;�s�Dah��3�Q1E�w$"5t��/��9Y!��Ε^V\�uO?�����Pl��^R���"]#�'��A�a����;�-,���O,�o�-�$qJ�а����l����V�@���h/��G�bxM�: ˋCM�z�5�%E4y����@d��)�h��da2�(��D��D��3��>���(�`q����]�K�E��m��6���J�JB��$Q"p���2x��	���2�H����M��ͱ�&�d�����)D�6v܎>!�3�(A��e���/��uc녜H�T\��L@MV�h��#9�}������S���|g����An��ڱ��W��_k���pw��"��ea|��~KFz�[�Ў^�lj�����b���;�w��"��XT�G-���b�j���ɼ�I��}�dm��A]�v����0���B��P�fO;�.���G�w�Nc��a[K�wL��э]��։	� �5u�(���2�������p�n��ҧB��;���\��Q��t�|����1m��~���G�絔��L0�&%H���SJ��=19h#PMN�򓊂���-#��/�"���哾��Z.?s�f϶y����n�L�?���11н���Y��XZfi�3�XJ��ES�3����h��dh��1���� �MD�9�S�$�Y��L���<��bLE_�e����8���z�>��)�q�A��z��ӊ��"���lVŠ��g��A���
/�m�kم^�u"�?+h0��X���3������x��?�OQ3�
s����&�g�9�w�{5v��o���N�gU���W QI}�	�	XLCU�t�@A�D'fg�:�)P��=�?��ƌ���G�9L��edҮw�?f��_��5��k`DT�Ђ����� @�*��d�oMR�)>�m�6�j�֣M[�[�����eB�'�����_sgģm���r�F�]
F�_-��5�J�*//��'!Mj߅j��5]BY�G����.�>]]�]Fw�a�D67?A�-���HI�ق���fȵ������J��0���E���`*�.dv�(.�WWu)xR�Ru��J7��\�O�р�&D��%�2F
�ī%�zd���� i�~+y�C�^�yc��'�ܶ���U����mI}:ҹo$u]iDz}Y���8hQ X�����b)䂜 �[� v��#�`����U		�x�I���=W���{WG��VIG^W�*:h�%�;6	�ՇҠB��$���%J.�P	eK���gѲ~���$��߮��2ٜ�]��)f�F�*��3ɣ2L6$�ɼ�挧��G��]#�N�~�t����!�Њr��	�&n+�ȍ0��dT��Ñ�XI�M���o�Џ���ULa�\sg1�G4<<����9V���]A-��L�~����s�(���:��qƏu[�ѓ �)����~����dj��P�m-�9G#�Y���<�r����if�K�Ԑ;���>����.#Ai���\����)Õ���F�l��G����r�j��h�*/�6�}����h�{D�v����2$���xRn�493���U�;�h+������8���u�!��?�
Ģ��^@��[�%CZ��-�@~�"��2�΄��/��JL�ʗ�ˆI����/[�N6�S@�R��>1&�#1l�	`A���� @��I��p����?�@�̻�ڦ�)W?�uc#�S�
�'J�3��=����b�Łc���*/��l�ބ39u|?��2Q��3�d����;)K������e�-mcT��^��
��z��&Yrr��h�C�̣i��~3�5�xI��!�]�K���j��xpp��%/�g z�@riCi��!jR��%�V@���x(m��-��	:�Q�����iG��h�˾��E�߷l_{�hضX�8���^�5����B==EY��㕠s��sU�O��z�9!�4�t�\xt(>	��`8�\�����$V�e�K��g�B�- ,��v���{N���w1��xF'�Z�����镾GM��dW|��A+�v!
��jO7��5[I��/�f)��T#O�su`_�}����ϙ�F�'��&b�.��b�������{mB���+V���3�W�YD���$�e}��o�1���{fI�ߥ�]lͧ�c�p����JH��U��F��Z@p��[2������$��\��/r�-���A'�)x�+g�#�3�LqV�a����Զw0!�l�Q;�uU7C����UG��ɔ�!mzr�x���$=h��6�ۜ��`fv
_h�F �Y��;O;��_�D/`ZOe�'(iS�N�����9n�ft��K+��6?AY�F ޅ���.��T�;;��7��S��y��?=�_�ݘꋡ^��NZ���6ĭ�~�=3O�38??�W�] ��q�@���A���G���?}Hn�3?��GZL5�޾E!�J	n9��څ���'�%+�\���6޾~]3�uצ��]f5��ϜShjh;�w��P`RY�1��E��M�|���Ґ> "�@�i��(����?�o{QfY��#��Q��O&�	+(Kx�c���	9>�P���mqi��x>�n_�^�cEn�+�&�n���gWr/�{���r�V��oѐI��ԓ"b=����6�� 	-�����C���$����ZȾ9��������&���;��}�˳+���1�oh�U��K>	X�|-�d7
�����"PXQ�|���*M��Zv�[�#U(P]*�7'�"ֈYPǘYㆻ��s),���=��n)�}6�bTŸ�F�=�av؝�	Fq��LVF�ӶfP���v�k�z���:+���(�<�.�Q$�a�����L���h3�·'��[����YVo��x�w^�f��6�>���'2�iib�Hg�R�+�hqGD���f^�W	J��|��%pm��3���;5*#C^8$G�.�>�3Ɯd�|����!j�l�y&�l��Hɶ�dhAʺ�-��4�H��z!<�4�io!��I���z]=`q�|�$�tۦ�=��>o�5��(���}�RQ��� |���s��Z����mC��J�X�˙��H�,+��+�ìou%��)����ӓ��<�ͷ>5`�l�y��� } W�?+�������x�B�7�?;Tҟ�<�B�X�ka$���D1��%���=��?�(3��&��o�ZZ�mW����>wo_FAW��s�ؔ��`n'B����5`�,�=��Λ��F��BOY�5���\�C����N�e�����)��vV'bh��s�9{5!�9����~An���#�h��{ 82���wțt��y�?4�*I��_�0�����M��i���4�O�FT�D, Mc�+M(��C�# ϸ��h�L

�������(5�G24�ې�</��*�l:�`ARz@dmM��@����]oK�<V��S�H�J��^+lnV���ln�K�}�=kܛ ����Z�@�:A}�}e��#��n�Q�Dc_��bYEDX!P8�j�����[!b``J_�3X���g�#\h'�}g�a��p�W:^m�/�� e���x�c��?�l���K�c�g'�/�fF��� �xt�"��J��>Q�!|���*����nYǴ�$?���,�n]����|�/O?�Z:$���\	�/;�5Өm�w!|[�rTw�,��[P@� Hh���o
�V0�5�GFD��%]���w�E�^�y������gN$D�R#{��#� ;��,70���&Ch=�W�s��C�v���I<��J���­(�D�\�ᮺ�6�q���g��v��=X��B���1��������jCJ<sB_[�V$:��S -�-a���쑆��7F>m�?F��d�K7���R��뽎V
K,3�ūK��S(�{��u/8���!�g�A��cq������A�����QG#G�X>MMe�H-M�o�6l�%%�������"C�:k��t�q�U�������}�77�N��C����U�U.�5Ȥ	�2�J'��n�3x��0�F���`s@���3|Fz�2E�]Y�h;R�b�"r�Vs�n�{�O��~���|������S�MY�����:�3����n".�@|�f�g�s�%B�
|�m/C��u?.ҋ\L����W���^G�u��a�퐆�Y���a�Z�W���S2+x�����`	V�?C�U� �v��6�0��h��by.�c0�!"���<2�����"}'*P�z�#W��s@~sP�/�e�(�J�i�e.iC�FQcf�<��$K�tgr���h(���J���
�Ue�ɨ-��[��V�[�����z�(7�F�T��{?�����ښ�CH�������)@@�oT.= �s��/����:��E������!B#��j0o�J_X�����ǵ��Lh�;	k]^��g1�'u������$i������l�l*!��T��#p��\���;�����V5pH:�W�x^5�4-��ޞ'�k��r>�vP���ڐ�I~ItN�Ed�O�O�%��L>���J#NXq�ĉ��|�RU�HG)��h� ��!�]�q�Y�Z�R/�����g�����is��3�Ty�&��@� =�n~���#�z*^��D�xte"���
�𽛀L��P' �Q&,'��J��P}?��	��N�z*��֬N�/z�8�% 3|5�������.1ջ�S�P���=1���F�;��"w�ѣ` H|!@~���,�ʰ�?m��xS
htb-w$I �ޒ���0�#I���x6G1 ����
�~9'�5��M��� �)�9��+1��1A��T�s���v��CWf65���bc/wؔW�H��z $L�}'ly� ��E���)���%�KH�!�s&E��C����'�>�#/}��7�3�SN�%�	[M�?�θ.�7�Z����oXX98DC:��� CV��k�?	�"I�M�%t+Y�x�Ǒ���t�c��?@���79���+~ ql��F��\A�<l���g�uAXp4�	�Yc�3�y�*�)��T��qj90)� �uzS�����"!&(�'�ux�
��%7��e�m٢Z�E���(F��.��Ƨɾ��3�[rѨ"@��M}�җt��?�6�&���zy����V�(���h{Ե�Z X�Stq�5��$ �ܒ~󩨮k=6�6��XF�j�L���:.L5��5�̡Be#�w���Jo���_.70���ݲ�Y�y3�U�����W3�n�y��S�7�\p�'bcc̓���&����h}_4�N�S��TB���df|N�4\�՚P������c�1�q���� F�]��?�ڎ�sx�7���Z6������U�Z�Iറ�D�h��H�Ӧ�u�%�I���o��l�>(�m�pؗm�����Ϭ*�t�p�ߌW�x��"���֖*��	�����8F֬Gl�Q��M�?T�Nd�	ډ���1T�xj5$t��U����Z��S�xf��݆o�F�w,�9SdiЄͯ��t�3�M��8��H͖'��qβ�"m�}Q�d�?�N	��yT���J��ttt�kǺ�lѾ2ZϥH�:�Wk�$�h�>�(-� SQr�5Q�����G�Ҡ'ǯqW�Y���^�O�CE��Y�`��3l��g%���\���Hw٘"�~s)�?�
<����Xf�1��1䦷�a�n��z��Xr���de�%R��b��I�����,�ж.1{H$�
� 4�+� YS�+\R�8�*T �i�ۅ4�}�d��x�Bc�gJ��*�6�����G��ͬ�%wɮ��^���1�OU���uK��P5�ZRs%�}*+Ұ��N�R������Pf��  �<�����˓r+�΁��`���š�7� 8�=U�B�D ��{}��V��5X�޼�`�刦e�=vzw��>�� �VΌe��;��x��o�Q���ߥ%�VJ����.t��'���"32�h/���}=֊⡲�tϮ8��0������ x��gG�~��j�B-Vs@q�JP�w54ygd1%�X<�&�X2C�-�"���	Jh��2�]�&�MA����z��AS����A��~��r����A�p5F>��	���RR>�/0q����|y��#�N{��쫨zR4��.X��p���<�����kv=��'ν$?P��X��4��iR�rC���0n�)���W��K"s�4�����G���,�^�!����]���X`�)�����cV~"��zۥ�a�:F+	Dn�Eds��j.WJ9��g.?�w��7�V��F�?�Jwy��!Ջ��S����&��D�׈��?
-ȑt�[G�ʡ��ʣ�@�_���O6�u���g��n�;,e8�vu�zsP�Irf�P�5�~���6�o1etf��߾���C%{��zeZ+g
3���C�pv��T����.��5׮oȶk�B�B�X���6b�Ҫ�=nx�3I�5�^�[�
n^��s
X��}'��);���#�`yTM{�A�>'��)F=k͎�bJ⥘5�b����Ț�����N1S�)y���������5�#��<o��	�����			M`�o_�ka���sb�?���6^��ar�!Z��PY�������l㱀#�g���;���C��A������{�f.'8J�7�<�2<cY�8DJc�2��I��&�ڨ<������i00��[ qC��)񯲨�ݤ�O}�����|E/ �28��ָ!�&=�s+���C%P%�K��Q�I��t�iM{Ğ�CD�Y�v�q4/��q�4IaNV9E/���eC�Xb�w�����e�m`�y��2M���sH>X}�.䤀�>5e��C�3	��C�n�aB�	{#�Gh��0(����ђ���u�u�Lx-:������sD�"j��GN2CY��Ce�7�44?B�>��$������߁���0�s�3�ȦVݔ 8GOՉ���'�F�91U�9,#�Ǫ��Pl��$�@>����|=v�Ҭ�X�p�~���ѝ�u�J�wtp ��r3�-^���{`��9������=r�����`� ��9�۔x$F8�j���#��UB�"oH��ydC
_��:)rAV�g��Kyj���Ǔ�;�)í����B�d�Q�0I����/F.I������t02zj�~h`�?[+�=�L��&tr.�DB#b�)i�д��a�^X�6�:Z�(Zz8��9O���S�zz��m+]�.l$�<?K���y����ei��Sx�_j*�)/*Gw��mTF� ��}��88[�7��L���
);̭ȣ_� �_�Ȏ�*(a�S(�{��';	q��٩^�۱������5�rDw�y��4��_{�E�D�E
�6��ÿ��m��KQW>0*�������8�a��^o]JO�;��1V���9T�����\�ü�&'�.���Do8�K�r�YB�;A�^+ۮ&�4�A�"��VM3Ĺ��. ��G�`y����$w��vܛ91I�gϺ8#��  K�k*�lBĺF���P,�Im���C%��
%�ٍ���(zX�b6���Ʉ�Et��&���|�_.�]f���%Kw~��� QN�	RZ�,)9����� ���p�M>ۈ�h�#=̿���q0���^��K���v��?��q�iɺUb��'?�O��x��z�����r�Tf�#Te�kD/�%��Օ,��P:�������u#���	�������y�1+D��yn}�c�V%nv�� ����j�����LM��.w�6w���3��b�u�6�n;��Kq��a�`��\�+�1a�3~&'��S�5�������Y8���x�)���FK`ﬦ�&��Z� �}�nvF|���IWp���'�Ym>�>��5T{�5���%���7m���������߯� �IB6L��b��9+�i:{}�d���-#�^���RJԫ���7	��bz�F9�R�A���<;��e1�q��М\��a=x)4���h��.�M}ц6���V�!�םSiE>�g�SJ�}��!�V��u6@b|���X��~�~l,�/xTQ�oqA�@O�ґ�|��n)�5ֹPk����%�=� ���ta��8�c� ���5/����e� ��=���	�����f�����:l�&�a���AºqblPC������?����KW{�	C�|�YL��Fh=L�Έ�uCv_`���~ >LDL�3�G3�*vNhQ�ɜ&�ŧ>�	��0[,ߎC��	�3�X�d��T��h�3�F����EH�G�˘q����d1ˈ�Ӆ_�}�iq�D�XPpQ�9���C�b;<������Lg�8�]'��4胃�X���`����)�5��Jk��z�L[�^_. �������x)�`�������N&tC��R��WOp�A�2�~{�if���2��wA{(��G�E�9/mptwΜe7zaT	���Q������h�qT8f���i�
E6���*����_��P���7ڶ���\ǮmJ�c(�"��F@f��KDf�sƗ����Z��v�[�l@]��	8�Rҁ�;�4�H�t&��y�`�&�&��[��.ә(�Ie�~��!"5���>x������$�0gj��g�ҵ�O(�fv�)
���gz�	�m�����ǩ��Ju��?�F����I�
�1Fk�ݳ6��f���^����:K��c��rk��wNK����쎂cߧ��ƻNЖ�h�}�v�!>��MM/?�~�(��s]bޓ�d��m#�8I��m ��|e�����E5�B�E?�/{`��V�eY�!OEV�c��a���{rc!�3����	�>� M {MC�9��2D����<��g�������0Ǔ�p�|_xA�=A�V�;����{8��IA,7X�*����������hRb��3vT�b|�;�U���00�c��\�@�G�>9�?�F{05����A(�
�L�j�}�q��v�lmx�&W�Et_)�L�T7�|@�����D���9kt�Y�ߧ����){�i�[��&>> �Vx��lk囃�H;*{�,+�|�5A���Ok������@JFy�7�5���C�9a5gn��T�!`E�U�<�>���AgB��|�[�nD�EV�� ���O	������t%����+�-�p�1������rqZ�(�Fإ㽐�σ�
C Ϲ��[�v)��X� �9~�}='�t�Y�n����]|E��ޡ�}s�ٳ<dI��K*)�.�4��\�!"@�����P��T](ҕ�FqG ����w�qp�o��Ԭ|����m$s�Nz�tKj/��JXE.z� h�`큚�w������?M��N6^��t��	���R�/�MYx�����]���P�k\�I��|�Q�K��G#������O�2�쀻�ν����SE���m�|��9S_�·�9�xw'�W{Σq�I��:�F�>j��W/=v)�g�)9ԠM��������ĸ��G���h�U#�@�f�����)�q"��UՇ�9(+g�\g��[�*g|�� G�e��'g��fo�#ʔU\��s��| �Jc���8W���˷�2�� �$g�t��<agY������%���틋�֍UU��/�����	����jr�����/b�����`ݽr��sUcTq���rY�o��[^�E��N�O'���-W��|��X�٬��wy�ݢ��h�/��A�@`��I��������9�����<U�^��m���n�z���Đay�����>����Ѵ��.�������a�g���[�����&�g1;N�Y�`��9���PI�k�Z[P�r�r�ڿs� A8�k��|� �ā ��MWN�n���Ppw��f��J��
�G�3���O"�#��M�|��J��݌�;��p�6�Op��&���j}}�$A$}�N@_v؅?��s�����c� �H�4Ot4RSC�|�
C
��B�{F39����w�H�Y��
��#������nYu�Ѐ�ܯ_��������Q�\!�;���%��K6CB�h�8�zZ��?b�������R�?3� ��k������4JQ��FV��3(��d'w����j�{��R��S�J����W�TyC��U��F�E�mo�%r���-pV���.>7d�\��������.�ӆG��[��
��OAK^�*�b�R�����f��sܺ�S�ч1��Z���٩:@�	�V�����$��1F�G��,"��x�q �a���M�6��0��/��5t{-@�v���`/�b�����8
_y[��a5��k
����-e� C������ǖ+���J݈d�J5�aU���Dɓ�M�/>]):wn��	�"H��03�&e�5�h��L�-]g�.|������5��^���.�c�����X�����:�� ��=�q�k�UI�#�߈U�U� ��}M0ѻ�kM��q~{��쌞g_��iî5�6&� ǌ�}C��f�vs?C � �"G�� D�X�Y��,LZ�%��y��w�8���&j����
����x�ʊ�P��?��s��������vӋX�M'Ϗv��B�v����H�ey΋���&���?Q��Ԙ�p�A"�F �?X�+hL1rI�?ҐVg�D� n[Њ_2���v��}�u���fJ�b��G���<�;�&i��|�6 qƥg�k/_{E}6aY�0,��m��>"F�@o3�s����\�(.�n���][뙕�a�{�=<%7jý9�:/'�ƔOC~Wձ<IS�
p�٘�lV�����_
�򀿙�/�h�L�������[�����EaK������f�m��\�t:(�
�bR���z�
ƅ��ݺ*2�7�u�� �gѷ�HSߒ4����o����/���|yM�_ �	L�/��z6S9	D`�m�Ň�o���&�S��C"���8�n���U%�U���L����Z���M�\Y_�7H�!�Ms)��< �/�� �C0˦_:��8E;�����5������7�YĞ3y�}��zwT��Ds;X�zHq%X��$t���t�3�-8�F�묘��� ������X��-Ib@�t��%��TXC�P� �;?=�22�
�t��q�gjX̙�I�|ڑۄ1����UdO��H�(�e��dÂƲW���ϧ��}�a�Q��_��Q���U̾��^�L�V�D�Mp'~�Ԅ~ �����놳��T��h�Q��An��=�6�l��(h������*�	�@����"�N��a�����wqOo��Wɣc�`������}O(�p�=��J
���wn+�W���mW�vI��p_���R�%f�hD��E�n��!^ n����){�o[���5���	9������������FΊj��g�S�X��Hn �ܟ�����Ak�Aϋ�����J�B�ŏ �C�L(�u���_f�m嫇[Y%�uqC�h��
���A�r#���	����S�Sn� �Y�v>78��oO��0:t���5��&�~9=��J�,m�1t��f��P�P�/�����߫���G�"H)�4д1��2_�.�޳��Nl���K�����Sf7�S�|��N%sy�j�> �z)J�G�@���]��/&<�Cr.��ͻ�g� �To&(�#]�}�.��Nݛ��2��I�& �f��}"!6/aZ��x�)+t��RX��$1ǳ�kURTr���_l�a�;��[�͟�N���E$�7D�_�{Q�#Y���.��*����
+;�"����d�M1V��	V�|���!?�!�=�s���I��]�G��� �e��	WW�UZ�g3��/<�|
�L�n�Tm���$K�026��� ���m��{��P��0p������m#����ӡ�B�J�03����b���a|O����7�=B#Ytрh�#�j�̈�n�?R"���#<��i��z@��� �M�
�S�-���Z���% "�n������-w�+i[�^8���ܸ�C�����|�}%�f�6���hB?h��#����e��^7�MD�9��C
f<��p�u*�����j��^���K��lt��(�3n����uC���F�[?>=0B��҅Z)�0�j�Rfu��z�,���>=(�u�%�g�Äz�������Yrю���+CZз�ϒ�k~Mc���ꗌ�����o��a�^n��x���F�R>#��=�V�����F�J��9q��dW�̖�+�;.~E�m�taA�6]VYTY�p���񃽭_1,�|%�CQ�0��''�ʲ\�+&6|N*��U:���p��w�+G�`y�������I�!�҅�+�0=��;83��Cq���Uγ��
o�g�*�}���l��L�U�����=<Q(��(>qt{lv����F�a�W��mn��v��^���%{x{�D��c�:��=~�4   ��js��W������>̄�"w ���=U�-5�N"9���hd�7���BF�OTR�ϔʏ7NF�d�&��-s�#Ciۙ�[Ӓ߳M�(:���M�}��^���?H@�}f�ܤB�Sz~J��G�k�"G��U�=$�.�'r��k�N��%�ڽ���|{�G+��qOٯ��x�@Kg�!�+�8`wvQ��0
�uJސy]B*4�QT��:G9E���t��hzM�@�'d0�Wl��"riX_��v#��+��FF��3˳�������̦sнA�"$�"�ŧ6�� �����u�3J}���0���ה?�Z_9Eغ��q����G���M���>��d�)��K1j�'�������[�;���p0&���f��W����-��=�h�U�������W�`����k���1Y��nO+�g�Z��t���0Cr'!d��%�v͔���:R��
X��K�Q���to=���]���E��ź��w��d��Y��J�{�Cϫ���S,W���\~B6�ѧZ�Ĵވ�YK������G='�����C~���D ��łl���K�Hݣ�|���d�L�p+��߃���|���8#���}��6��Kţ�R�!�}	�'N�`G
�sA�|�:n�@��_w�?0��{n� %���A%��];V���^�A��$s�	�U�oƕ̪`T�c���s�]�����(Ǥ@�Z�ˢa���NdN�z��bt%�l�!R����0�{���AN �W��n&����ߚ�l�_�M�]���pk��+2G|ێSds��\��n��/�z[���^�]Q��1�!4h��5��8�S鳙*�#'!s��RB����t.�{�Q���w�N�_YY��j�`0 ��A��\��j���]I&�5�\m+��(��6���Nvl�=������)�z�5������:R:<9t5���-ϋ�kY]F�q�X��:��=�³#̤L� �	ڙ{���ivӚb�1B^ȓy�sړc�4�+T@�ႆ���yT�-x}c#�˳�  	�N��Y�C��K��zO�Q�C��hۮ ���A.����w���č��I"V9U�;��p�������oZ�|yB���VyR��� �G=E61F�5�尷�aa����1����ƿn�?������,��蛺}�E�� 9�\�KJ�B��'�b]ؒvlPy&�L������R��0J����s3վi��e�oWc^��Sd'C�Ռ�4����4@��,�+i<������Q���s0/��	:���~��O�;7���c0kV]}%e#��g�}F��Yo����[L�Z�3�r�_�<�3� �dѧ��<1��+$B�)�7E7;�b�U�զ,{O����&��-�N�2�+9��uwD"�X�L�T���FZ5�Vk��Hh4"a=s}Wd+��&4x" j�V~`wx�n����0qm�>��s_%���Ӻyt��)E?VW#)[��b�ЄQ�;Z�����k�i���l���ܹ���l��L�Lv������YLPO��v����k0��=�=��/B
S����J"���0w�S�؆��qB㇀2�F>����ړ�Y!�r��T��@�A�Q5��8�Y��������P���x�q��a��'%���9��W:z��/��{}7� �.�Xwh�58앥A1�R��{�t�{�U�r�J�/��p��z˰8�%Zx�`ap��0��<�� ��w�������;\r����}���;ϼ�]U]�Wu�w&���e~'E/D�s-m���a���_W�(@��s�`�����$U�bh&��So�����S����������Ԫm40'ά��7���K�ơ3<�1wA�%^VU�z�.��@�҉�#�y��J$�_ԫ���%MyyjQ97�h��s넇���ۑ���T��q��|ľy)��)�����5���S�������w�S<���T�_Cc�؎���DU���s1/�p�<ha��e�\�7?��K!�|V������H��b�y5eT��sA��q��e���h�.y���S; �?����v<jz���nHZj��\�DL���c◄{�z2��f�������'�]��<�:.g?t繒Q��6C,���܂�*������[pYA����Q�eG���,�c���_h$�KK*djQC'�4��e���v���o�������N���Q�豍�����vြk;�:
ˤ��}��ٔ/9Q�X]���|
1hRBA
��l���&*R�>�ll(�_�Any(v�]���R��Ws%��-��н
�7{jR��������7��e	�.���)�����w�
����e�Lu+Q/EN�~��f���;f��d��n�x+Y��R��O4#͔O�/C��O$�"��-��p�����=�8���B�	=��ǫKI+[�,��*Z�Q�a��]p�S�F�T��=�%��(�o@G �)1�Kp�j8fp��ol�W���IϑV/��̕w��蓔�4%�P�0���%Һ��:oR#Ƚ�U"j)j�\���"O�'�r ��p��B#(��E}6�����o� 6�MV�BK��M�qUrY���Qy" ����Z��������&fso���ň���i_uZCa�@/�58b0l���XeL7��m0�iJ��.�$%�[sOں&��/e�I�������~�u��(&�w^8s '����
Ę'��<���t�̹�2Ms��x��
�/����~	��D ��=�ψ�owUU�F
������HCg!����)O�?�9ϐx���]�W+R���I/NA�������ϼ���㫗r��ɮ�jr=���2#���~�j�ǼbkP�뱦��]������6xHQ}ة!?!H��ؠ���^����.�T���z!�S/6q��%�/[ �K'�.I�P*� E��{Z2��qH��7��+n���osy�;f&��W���h��Ġ0�κ�6z����ދu�?�rU�3s�P=�w�Z?g|6�xAb�sZ�V����<ɱq�7h�צRY�8�_M�8
*]�o~D�?�-&���M�+���B�tO��a>e]�Ab�_EM�~��A�7�)�N�/+
��?����]c��5E`}^88�0�Xg���]="h�L�1l�X]Z\�z\�k�c��ET�$�&���׬Ԧ$="���.��қ.8��M��M�Y\�Q�% �4�^���:姼L�z=�Y9ߎDRKqә(����%��'_']��4�H��1�y��¸���;:��-\�����j#��I>%ҋui(Ok�5�8A���%8��1����t;\�)+gű��F������˘�w����&�xo)�P-"��\ݮ�w}�N.��WᎦ�O�_;��%�3 ��m1fjvػ�	8��Ji��\�I<>J\t=���jY��[f4V3r��H����^r8Ӟ�_��+����w���Zl��8��C$$!@�|-5ȍR��2SC��}/�t1��~F!�N��KF�B�L�Q��@_�턔�w��#�D����Fڠ��I�r��6�>�6Sy�����
�멌���3�A
�̪�)��bdf��Ј�@}�3	��� �}�X����Z��/�w�.,r�s:Y�;��z�v]R<O��rW_��D�����^Olʞ����`��z�a�E�}�۹�d��R��}�x�iN�3�	ս\���1����������}	�t񼄴˟���c����!�;[�,/I�m��k��Bg1����;�TpE���a�mL��-��Oط[^��?�zY�!bVΗ������c*#���l�~	G���2,BU��Zn�^C��b��pq6�ud��
�W_ͽ�s?KؔԂ�z*(�aS���F|�>���=Y]��r >�{��cj�Y�M��\�8�ZD�tE+��T�C�s�3���ڒN3�����i�����Ĝ+s�/_��u�?1��S�z�%Ӫ������v�_��LG�B�5���bĪW�;�)K@b�\gh֮�z�����@���D{�B��Õ8�#���ϝߦ>�G�1ʣ��[�!�v��զ��r HB5B�ݮ�)��
A��a�;S�7N�[�V���{��t�oq�9�����l���}֑�v�����9]L}�A�0T�E�����;Cj��
E����	�臿�m}!�!=���	1����e����1P�){a��qj��Mk���b���*�
���UW<8���KB1ȑp����o��x^��: S������\3�p���8�굇za4\�2��w;�B�����GY?K?k�s��6=�c�<��D�Ɇ�
U�D"�2�P���"��}����kݓi�@V�rJK�+���510�1�^pℳWXEaM;��iT6]fH��J��2*��GJQR%~<g
�q'���
���

��)�Gaֶ@9G!z�b�|ϡ9\��ۙӬz�wH�ǋ�0�����'ơ:ZD�͊�d� >�ޚX�R��OwY�`�!�FV^��T�iIh_����i�a�'�9kf�,��.L�O�Κ��eA�ez����S_�:�W�{���h5Ĳ*飯�!2�(|=$�yD3^!+��h��,H��S�	��B��>���,�y!IԔ7����ii{Լ��D�p�TQq��Qk�=�;��oR�r���"����N:�����{F�D��sl������U:��1&����̦�0�w�?����u����Zk!`�vq[ѧ����C�Tn�Fŵf�Bw�a@�*A}�����=	�}%.96�R���S�)�,�[k?\/['.R1�!��9_l��������=��ɬ���@�i�f%a���D%Ą�(ZQ�O���!��t֟��z�@�J/�� �������Y�b���HE�H�=+�X�~3ي}Ṋ����E�KÎ�ȑ��� 4�͓ScIa���J���T�Իܒ�F;u��Kwh��9���lqh9�phq��E,�"Y.b��V�/���4;��z��lT[�_ċD��C�>;���6ds�n�v�(;6k�.����Ծ�`fx�^�r��S3.o%n�%3�D��F<}��5,3v���Dm�Sw3�V�ײ��.�	�Ύy~�će~վ.Ar�=6�2�/�at`���\#x�w�接r��5�Ӫ��2�(G`zV:�1��}�&�l�{X�@��Pu�6���HW���?���|aX�b��}�}�	
�R-�'���u%:�ߧ�Ӈ}�)�&
�-p�"�8.���[B:��O��ӷ�.�FkN	!���ץd�;zM6�9Ϧ����PA}f�4L��eX:��T0�!�c���a��I��vV}`�d��|�D2P��-n�^���[;;ҩ����) 5F�K�s������Ր��2�4rq�B�@��'O~�e:#I�e�B�uPHn(�BfD�A:N2��;E!	��{���t�Ea;t2�E�$��i^O5��U�SL��.�z��8����)�����;���&�{/��.e��Gğ�� �S��F�)2�V���A�}ȼ�tʲ�R9�=U���q֥��p��������%ЗqD�n!��G���s�e�h���6%v�Z���_����q֌:�F(NM�O�J������N��t�:��?"Q�}��1+ %�,��q�ύl��ג�T������̊ ��H�NQ���o�'�:�F�ѿiB�Lw&��Ă�VQ�¹;y)��͏�./�{�/�&��������LQx�V�S�D�"��9�{x�*]X��n��Z�uE�1�����ў�����Y����$f�QjHc���P�9s��\՟X�o�3w�BJ1	$0��泭�^�<�*�r�;�5����u��lĒ~�Ǟ>�q��T�b2ձ�oJR1F�oB;)!��>�µ%a/���T3KaD�p~~C�;W[:��w���y�l��[^��Y��[�h3� �]z&������S��?�YD^���V\���TX�U�ڌ��媯qm/��e�=@�ci��R-�|�w47�:ϐ�δ�OS%~�LzIW˴#|��E��g���η��Wט�F�����#�d�O囹rA�=��ը��H^ (T�C�Ua�x�Ϥ`� �B��];�4D⤺��8o��/8� ��s8IN f;���|~ރ �Q���wE��rX�!#=��u�|h���c�|�T�r`-)��@$����y�L�$�[�0���*y�o�〼��Y�C�R3y��kX�`LL������x?0ĳ^����m�o�b�jQ���g��֏nc�}\gi���Q��o�$�[�
g�~�e�8Yw��p��}���j��.��D�/
Q�kB]4��%��%������Xw6�K,x���)V�1ͩ|�U�Ǽ����+a�[C��ֲ��P���J{�p�8���ե��M�@>?t��g��|zQM^8g�>�b�O!kaGcAZ��U����yC�w�����6�,�w4

��Pt�S����^�ε�rs�q�,;����6М�M$R}(y��4�{cj��j�+��oF`zjO7uܷ��5#M~�F���ּW���ũ;���t&J���4_cV�iq�0M���ɝT�ܯH|g� �i}�E���(�Ny�Lb��:�@]yc��̂�@���u��c���݇Z��p:�����1��p��@�<�)'�� 2����"�i���-Z�S\@�1�]
���כB1���-���eĺ<y�p�*)�f�T�|6(�URbMS=U	B�/�!B ]���@�E�}��C�,�~���b$��hو���_c7��)��|����o��ϯ�� E�?["�B�t��+�9K�D����#�^d��̈�_���)<�0d�J�rwJ�ـ�&��ln��*b����r]�L���+o���dcbw��ʠ�`�q+�Ud���!����y��B��^y����~��ï:E�Z��`eb"�V~�	����XWĂa�E�Wn@~�I�q�7~
��a"]�d��_&*'5uyUF^�Tw��ͳ�b�Z\F�Qg���a~6ev�_2� 66�bRv�F�<烅�s�C=�@���\PJ��H�;h��[����a���ԓ>�rq�W��?a(�ͦ��,M�#�Z���8Cp�M���o�(��*�Ӗ�^w��!��N���
��s���z�Is�G��ѫ�)/=��8���"���~k�_�o}��^#w}sM;��'@Ʌ�S%&'p���Z��t�2ݿ�$d( �2�p��|��o��┋�ČLUg�ӑ��	��4'���G�E:��0�.�~����M�aׯ���ީ����b�����"�\��oXH=�|����k0;rc��:s��)�Dw�zR	ǔ<�!�"�BJ|p.5��r(�-*���Ɔ�V��8���6����<W�X�HX�\�������a �B�^K���������g1�YK����>hj�6�ތW�l��_�iwJN�:H���v�y�F|�i(����]HއI��̶��[�P���i}����hZJ��_��jȥ������
+?ҷ�Ll.��=��~�y�Kҩcj�I~�܀ʡ����"�t/�����jm�������"_VV��z
V���󷦄r.������1�qEf���ʻ��S�^հ�܅�皲5BL4_��qd7��uE��7��S0s4�- ����0h$J�
�}�&��|� un �Go�8nfyc~Q���?G���O�1�\_&��zm��:0�;36^�R�/����̐$�h��I���K&Y;�y?fձ�}��7>��z��� �1Y��?�=�`��?>��3d�}� 
�٠4��Z� ���	��d�t},�QҔ���xF_a�� G)�"=���&��De�%����-��������7�\^^ ��,�2"����Z���,	y��4�C���ѯ�[��d��c�v9p�@�HO��IiU��}q��Fʕ,PP�%Z�h�4ͣ�Rc�O^�R �¤����r��(��e�G��\Y��4�yl8�Z��^F6��0�����\"2����WkAS���C�h
$�n��b1�/��}�v�"��j�WzK~Е\;�gș<���z��V8˧L��ܦ�>��Ǻf�`�>�FI��WH��(T.b�����#��Uսg�]pijCU
��: 9sꞀ����a8C�?4��lltx�C	�B��V��Q��r$IX
����O^�����MS~|t�i�9;����q0��|Y���NN����0����-�O�����:�Ag7��55Ԑ�)��D�h��m��j#��9�b�]9�/L1��_�6s���� vvv,Þ}Pͷ���_}�=&o�Ǟm��Ɗ<����~C3�l�{��Ԥ��j���y�W�_#.�(h��R;��Y��'����Zǂ����.CP�<���2�.�a?�l3�%:L����P�� ��.{�4c�C�Y	M��o��U$)�CFc�܂yI� )ق��ߏ�0p��O��jLB�?�V_&��{��*e�F�2����t�c{Ge��.dh *V.<j�hpX��x�KIZ��� �նH���(�r����<�e})k� �ҥ��"��c؜ׯ��U����'���7����M�Z$�s���c(�ľA��F>!�<��#�Ƕ��WUFS@ܗ{� �!uo��\�����)4��cPPR�z��9�&1^�X_F&@�:�C����yw8/�F�ON;�c��[���d���� �S�X�@����X"o_����
�>|zR[��iF�F�lZ��5I��P��ϩ��������f +_|����
6�H��-3d�.����G�f�f���)�41� �l�3���q7�E)1s�?vww�0�%/���% ��X��g#l��}r���JCy��������?�B���?|%g4�\(�ٱ�˘�h((+S, +�dYH��~��!�'V���g���
�`!cR����QC�mYA���C�T+@E�Z������1^,ݺ�!	ͬ��!����i�2Xd��ZnE՜����P�A��?�'|�So�h� �10�'����(x�կ#�J�>RЌ�麦��ר���g��ܨg?��	�&����PQ��I�z�k8) YT�g�k��q4��,��sf�'nL����\�o����?��R�Z�!��x��?��G���ˡW܊�,S|ۥ	��I��uIT�4ݩ�
A^"r�^���П�	��$�g����DMmv�����+1��oI���^P�"Ǿ(<^�G��!N��\O�����?�v\a�цg#�����RlA|�b��FP�����\�?|a�C~c�inO�G\�Vr�IlP��g�,�?}}-e
��D�mQKC�(~Ky�J)�	B`~���|A`��_3����~e��P�^���zꍐn�5��_$<�xjo�}��i%�_WZ_�ș�t�v:��kPC|��~thz�{�x�(Rm֓z����u�T�p��m�&Ri��t�db�k<��j���y����>2}�X���6�=�>ۈ`���1��W	 �>������������}򍒩���N6o�G	��'�\��kW�NrYD-/ԿpC�����>G��ʴ��_,҆�/G�@s�;�\�EsWw���L(�o<����t�L�<������)�������+c�n��3r�sr���$a^^H�MEm�0��^1�Ԣ&5��\�)V���Ρ,�~���թ4�^��('��]6��κ�����3�11�l%<Sغ`�J�u-v�RJ܏<�!���Օ�#S���m���O�r���>]�3�$$���Lj������u���Xݺ��@��D����AcF��3�-w�7/��c�yi��}�:{K����H��ǵSs.���..��Yx�R#���zDc��ޡ�|��(�[&~t�_�s����1�kn�1m���Ks������U�7K������6#�t���r�h.�q*_��n���!�$�|�\�ד����-��mmYĶՁ.����Z{5ߒ��/�`�������---}��iQfʒ�#�%�1~��N�2��X[�9������t`�+�n ��v�mi8I�^窽	���tF5���{�����0��Q�r׀)߆��nvĂzD~7��v��k�+�#C�ww�o�*�_Y Ȍ�Ͱ�hR�WTDO8o���vȨ3�m��Y���tA���&廄�K9ޟ������fc���.���M�"Ep����J�ǚ�_
�]7��k�Y�SC���Ұ� ��zu!�64��w��i�-����n�T��0ݞ!ݡ��x���q���[o���������� �¸�v���^p�����߿����!ٽ�<�+��Cy���D���`+�2+��#��K�y��}`)�M��I.���?���sK��H񩎌��x����MO������B�9��-#��۫�'�*�
��~�	��x*��c�Y��$�\l�Y�^��K�xhN�`pR�3K4=[�(*��7ڝ���>P/��Pڠ�{�6�Jʥ5�YM1ß��6��<�b���8�T�ڳƼ�o/WD��dN3�B�'�Eg2s�.'8��$���u��|��}���[Ȋ��5����A��40��>�XJ����%�u8�yG�{^*FT��3q�pQN7a�T��e�nT��B�5t`�ݣ�`xu&�!Қl�Lw3��l��ú&��.�j��>Θ���D�%;�W��;l���v��{8mV1�������{����H��~|#��+��B4��n��/���? 	�?5w���"�fz%�������_�´��{��F�^��z�5!~�2Ჲ��y�e�����Գ(���*�B���d�Ƴ-L럻M�����}��η:H��x)4�J��ަ[f�o�kV������Q&�]׏%r��	�\Z�;Z��ƹ]�ѿ�%Xnk��F]o��I�g!�ݲ����۝l^��T��t"�Z���_=��t���l��0CS�]��j؏�j�Dؠ�YB&BN�Ä���-J�?yb��2��	�tCMdN�@6ZX�%M���V�� 2z#U�����:��O�AR����K�$|����z�����^Q��ɇ�%��L�t�FD,K��ϩ����֙>g�gIM�R1�[�6�L�̓��j̆qLc�{|���1�r�_�z�Z~�El��_^��??-N�W�]����7j��t�u�����C�wu*��,��h����H��1#<<|kJF��������(~�����AE���H�������������|�ٮ����tM�3���ߟxͯ�c&Mi�U��A����5-+Z=����~4&s��<���uVu���]���{�ى�؆�[��dV�8ʝ����|��N���jT��f�3y�R>�5ʯ�v�(Gc�X@���}��m���m:�Mj��^T�ڏA-g�+��G���e$A;L�3	s�X�{��q�}9�e��~ǗΧmАC>x!���`�r�
sk��u/����ق9����I�����01��������Q���.z�0qq���Þ�e��I$�)$�^�iS�����Z$ϻ�1h4KX�:um�j��D����PM�P����� ÿCp{Y�_����{�>��~�E#������u������Us�a.b�&j�b��?,�����0F������~��1����N0����~��']��|�i7�=�(�eJ�����γn��?����v���C;e��U�8�m.ᥴ/������/c+H��:�?w&֎�R]T�����J��k�J�t[�֎�*�p3<rqBet��8�.���l$�o\����*u&I�n�g�"_�4}a�+ە��w)V��`W\w�3�]�!��S��Wz���=Y.{:L�7�f���x�v1R(����N�K��e�v�Mkj�Ϻ�:�_�)�˗F��/Ђ�=a>`�N���"ֲJ�v
K�H5GtY]��-&��\�ֱ�������p��bN8�����Q� �D�Q�f�ɨ��W�uZ"��è�/&ez�	�;�U��>�L&��>i�����00����y��$�ԕt�i~�;p�9J���{�Zbm���Q��w��jA���.��q���h��U��qOd�v3�K4�J�̖��9����'��Ar���뎓���"��	����%�d�
��ꕗ�z���S	�bE=?�<o��x���w,޷:f�A��?���s>��no�������*�M"/����a�=?���̿oʪm��ӹ��\�{,j����Oэb��G}|H����J�,:�5�_�w1�i4���v�}p��t-��ʸd!���JA� ����lP��h�t�~{�w��	�
6m�P��愁{��t��`qسu	�r0;<�`f
H<3�uu�h��8O��^�t]9�z��nˍz�S�>X�"��������*"��1���Fl>����O]�ݚ�ߧd��z��������hh���_�wՑ�F~:p]Nk^������b�ĕ޿�����b��og�fz?�"j�B�6�c�u+�z����z��3�נ��*C
�=6�9�����H巄�+�ʰA����w�y�#�$x�u;��`d��վ@����!vh#
m5f��I�}��n|�YȢ�R�+ao��j$�p�sG��"�C:������]������xQ�)��$�˴[��ߵs)��..��,E�3�'O����K�I�5;p�r�a�5'IZ#��Z׮�^�瘙,�z���}.�2��m_��G�[�<y��~׭}��4�uuk}��P����Y`[bIwkV�;��I�B�mFS�6�~n�Z�됅m�S�H ��n
@|ax�����7�	rƩ'�����}>/[��O�p�$^g�j<�(�a�C"D��O�>��{�.�Fȇ�4�Ŋ�ğ4�z-"���C��*�-�-������&��I�\�}����mY����{��9�ᒢ�R� �������ʝ�o�\�%���P���rS
�f>M8�}���W�BƧ�K�O[&�ҋ"Ϸ�k� ���Km}"`��iҩIn%����U*K��s��f�^v'���?�98b�y����kq��촉,?����i�tw�W��=��2g��K���Xz6�r?�RY���Q\�?��,�	�d��E�~���d�C�'q�_'I]��Y>o��75J��������%V���ױ��>cW�~[�̖mۛ�w��kj�c��/�+x4�X�(�]>����0-���1��q�g��3���Dӓj8"�����җ~K��:jڊ�S,�'��
�\Ԏ�i�?�x����#��,Q�<�,su��jc,��ޚ���zV��Ҕ*�s�	!��@��������" ��F���{�X��cB���)6�AI|�}�cy��u7��ج)~8�d-�)�K��Q�]7��۩;D^�LE[���)������jҿ�\�����X�횾�uO�o�np���/]c�"��W�Y����|������m�dg���>�Tk�
�o��="l�gJ4E:���ֿ��;��Vi7�'�$��riYw��b���&�R��N���Odܓ���a�@7�XJ�T���_�?>3D��O-uh��{�Ð�hJ_3A��?^������iX �ٺ���)(�-R��Б���oe񐉖���ʯ�Z�N�Z���F�X^�D^�*΂�>���>Ȯ���~im6F�͂%����U��mp�9��ܚ��L-]N�L^�ݕ`�=�����OQ�h�#ɬ��Di#]g����4����'���R04�[�i_�g���:�L�l���~�YD��V锩�Ǻi�I��N_���$��H8��z�3Ru���YCi�X��-#ǀitE�Z�-��zw�7���ҕ�Ϥ��SO�)�L�uS6e@���3����~�e$���H�i�&�Dz�@ϼJ�=����fcf�[lC"mPΥ�nW���
�Β��߶���Y��,j)�����οS�0j,���L`a�}�T�%	#A�9��I1��ć-�Y^�q\���io;{1+Q5\�0���)��F�ո©���N2�����-�l^��f��8�ч�Ym���Zz�$T[�~�U����ſ�˙�9�0A�bbr�mKW�f�4A�����f}���1��^ăV��,I�_����ҩ��ow��6Y�����.���wE�/t������X:⧂�#�,�"9O��$O����L�k��Z�8����.���i�ħ����Y1���y3�㴰2�((D'�莚�\�$r:D&oߠ���je�6�۪p���.��b���ܫ�iȞ�̀��|���fgoK��Mj��m
	���W���WTB*�6��
���%��,�
��Q��*�NȘ:��C�������R�ģM�w�� ThaCF�=_��E'B����B�Z1��TuN�����U'Cb�,tg���*:C�V���x�O�v�R�b�a�W���m���Z�������cZ}���GаAib;u�*N�tR�壦�Jr榅(���l�� ,d���W��eU��A�w��gO�C2�xr[nA&�/-`%N�<\V����S#��)� ��`=��j���������-��ɷ��$�<}T�G��䘉����!Ďz0��.�H�Ɓ���2Ky�o��sУ���f��-'iV�C�l��SW��O�r��"*9�����D�
*��ԥ?�/�g'�-f�-�4>�2���y�����s22#�?L��
~�l�r���������w��"4�/Vj[���E٢�Gy��,Bm�2Y��Ã�d�Wh�޹�Xɩ:�Ҕ�`��{SIJ0ai�l�����]�#�����Q0��( ؉�-�{w�Hc����cʾ�[z�?���k���y���C>?οK�NE���S3�FƜ�2��������N��c��pl����D/`^d����F�ۉ�&�mٺJϷՒC_R�`^\ס��hC����(��}�,�2�`D��c��������i/����}:�$O���<�b��H��V��'᪑���r?n�Ji�,�T�������?uڙeᱫ��MD�a:����>��t�$���H��y|IfI�u��w�ST��|R,{8n����3�k
AC��Fs��U�g�_����L�D�:�O[`	Uz���#����"�Qh��LA
G��fu���R\�616`LgD��vҾ̻�CZbs��TБ�� ���ԣ�H��<�6IO�����2��1��ULb�|x)����Z@����h��#u����ڱ*̰7<[�ݡ�PIݗ�ܜ��+���M�rZ��^o��\D� �S��Q-e `�h^��w&�<gHس�i�JD�El�z����x�H��~��??��J��3*�t�����D6�؆���wM�u��Nn㫌̈́G#R'Q`���]�!��5޷?��t�4֛[��s�4��7ŝ]�M�uJ��N�Y~r�7�M/ͽ�3�M*����&;��co�9_��g���gĸۥ3o��A����?����FǓ�X�Jb9�7M��O+�`���F�[N (��r�/q�'<�JmX,�xmZyj�'�TA����g\���������O���>l���@��=������PK?~�o;6h\���FO��"d��>��t���i��֪���-���<�o�����P� ��I҈�Җ��ck�}�]�t���1���|����nf����<�g7�
/)K��}1�v���;<���4�D��^��.?7���f��'.��T ���BR�6
q6�Z���|_h�o�)��&ə!���tt�^Nu�n�W��I��]�����,�>����΅J��u�w���O����O���o��cE+(�w�&}i�yggT�1��g���L��r���:[T6�j�u�����rV尠e�{Ά,&�?��4�ٕ@^�!!��ȩ��h��/g���{�q�ܠ��i7��R��7��C�RM+��ɼgµվ����ч�z�n<Wnu8i��\G��C���EH��$���k��!uW�Ta���H唹��\ܠ����~�A~���0��$�����n�{�!���*̅i!�J9��fq�6��7y�K&�	�7������Y8]P�\^�;jo�2�9�\���j!Ỷ9y�E>\���P�Ʋ1��n*޲w�砢��B{�d�Z�f�į��{��G�e����l�$'��<`�f���l� ˟vM+�r�5�����پWرd�O��&s<k>�l�c�Ov5?�Ij(Р��� ��y�����	�q*�U�m��82B�,�z��}�<�c�+��ܓ�պ�v�+�tV���4Ő*F�W�_C��.]�=o?�����
B[�Mn�5\q׹��)�ZMst.41D�O�U/s�'%�K�c�or�r�ʤ�zݞ{�4{8͡��/%j	bV�#Op�R}r&�?O
� �ł�޶R�S@���K&h20 SFPt�Z�Τm�΄8��LM��>2���A��o*�MuI���e	�� 6n�f�̥f��g��1�{��P1v�m���*���z����`��G��Q㒽}��m�Z��A%�b��"jt�r��oW%��B�	���x���n�\x�Yo��D@�O��#b\��u�6Cm��ٌf}��iQ��eڀr-���פ�9�|gW&Zz�@���S#�>�z��l;�)&�����z��E�-��z02���*؍CV+׈��<no������z5����z��'�6���q���+�4���j�ƻ�=���$p����>x�u�7ڥ�h��D��Ng�L��$��;����Y�A��t��z1:I]}�5m�/b0��mڸ�ʗhL��-�8�o��O�&0�pkt[,(�J�e Ǹ�*3�{v���J��7�>zO/F�v��h����$�63��K��Fm�V��r}����������N{%��1��>Z98$�$�����8�&:䁞�N� Qd
QB,��ܟ�p�@o����e���x�.��{����]�-�����ݎ�Hl6�"_I������}����u9�X;l@C6�*/���щ�,�퐼�`�cd�D `�oJ���'r��F�~l��۾�QU-ҒFu�R����L����	ǔ��`ϸ6�	�Dݮ�1�5d�}�<,v�#$�:17#�e��Í����⏎�s�̻c_H��`L�C���:C�T������T��cV�(��j�j�%�5��W�g~ �I��])7�+�L�\y]���q��צ0���oexNܮ��\�׌�D[�r?a_�y=�آ9!Ɛ��6�*��\�+��7U���7���ՄNY�Ox�tWv�w~ef�{���<PD��/3�tem��D}("kݻ9�4lFg#.��r �'a,�ZHJ*�6�����gi4�[e�a�sߎt�^�����PsQ���Jv����{�񻌙
 ������Dc3*@��QX�����u#b��,#9�Q�����GK�W�^�~�.,Y~1I&L�g_C����e�Y&G�G���}*��0��j?r�k�\��t���e��8�v�R��{��+��*����6��]���U_�"7�< �7��~�d��y�K�&�f�T�`�n��/���ēћ�T�@	Cߜ������a����9=d���# Y]& ����mQ�%ڂ��S�c� 6�/�{��{	]Cgm1��c���B������d����4��Y���/�/�@�d���x�� (޴{�pM:k{��=��?:��1��O���j98"�s����;7��844���CQ�Me������+�%E�w��2�������$�d��5�D���F8N=�'��7��1px�T6e�Н�Cb�]Xd��q����R�\qDZ�G34�e���T$_J���-�?���!9��a䟀 H�𡖓c�>���/}lD<����mQ��9ā�/[�+p)��⽫,,g#EnXx�I	o����:����� ���x;>�E�GG�[���GCV�68h��P7��N�%�n���޿I{�B9� a�����pm
�ѐ��c,v0����Y�����g|���t�V֎Aw�E?q��5b.�=���ly��j}�Vggi<��0]O���G�G"X��:k^xϢ��������!\*��uw��bo'����'Ll������ �k���x�.z����âjߵa:��F��$D��ch���.i������.��CRZA�ށg���{�{�����5k�W��y�}���`L��V�i�a��(����_�K��������DǱ�se�_�(ԬM;O0��>"x���@���-VygM��=���?ͪ�cR
6��O�1ߜW�����	v��o�$� Ok~>�mM���\�^M+�
`���$6�rEq���Ug`��F���w�8�S���g#7��N�g����E�g�|�,��/��$�.R�	�c�"M��7X$#�/��A;k�O8��5��'���֏?�����:i�UX)0��R
1A�m(�����[0ɵ�"Np�8������\J>N�����ZO0��@�R�	t���-����56�F�kp��d�`���ԅF8GW� Jj�!�/'�B�E�h���>�y�� �H���q�P��Kq�p�Ȫ�_P k�3̧�i�,���L���O�v+�=��7�K֍�:�\�qK�k��)��T�t��"��b��v�V�jkhn\$OY������i5XiwF�%�H�ذ��_�3m��s-u������Qʪ%@k��P{��}�F��'
�Ҭ�'ӁCB�_��	�RIX�Io $-*��G��Y��<����M9�f!UA���0��c*��u�S��&���	���7��o��ͬ�i0��[�y��+h�a��p䎬���u�����qT2�%�ol	�bT8$G+��P~����D�X���%6�L�Ot�-�}����9-�������U���1�&���q��h������q���b���E&�Y��!���1A��Eɸ@��D�s�H�?H�i:G��}��ί��^Q;t�w.�s�V������f�H���z��Y�,,�����vw<ܫim��<�nexS���Y���%,tF���җ�{��{��,�k����:�s-hА��ܝ)�49��Q�n)���L�cL���L�;0���-���G`��
�۲O{��\�;b�����CF��Y4�ł���$x�È*G)�<E�%�脭>[�h�e�{�:��ϩF<�gU��ӬY�Y�:3J�\Œ<��O �g E�|���7���u�����1�N�OO����r�{����nY�'�͍�Dr�����QR���O���ɹC�|�D�V*�<�Y��ǵʨ\�Y�-����/�S�,�����-���EMT��a�$]tn<h047�c�&�1��hVbA�M����0��ĴZ�ظ�'�S�3���&�^����/(�2����� �M���<��9��v4]Շi3�h�*�<��L�j���-��W7H{ A�d���Oܝ�`��6�$�_�o	>�vq���hHYg�vd�M1�Ka�b�����ʙf��Ʉ?�t*�Xx����F�F��-�Lc]��I;F��x����aã[�����h���M�X�j�'����]bjlۙ?��ح�	F-�M�3����� �ֿ����Mvmq��!�ua{�� �d�Bi��@��.���YBn�l�&��ހoO��.s+F�����,�5<��r�
3����H���e��/���p�fI�{juV�%���������1�ƚR�ŏm
�ɍþ\,��2�r��a�$��> l\
�jA-óG�i��3:B�!��w���qV�D���/z����ϼ{g����R�����U�K���������R�
��?���4i*=d��on�ѹ�y?�'�3.ƭwY[�+�>����e�Nn��no���4�������c,�����X��:�������8������	�*���pr�+�+W,�*i��� u*��S��ճ�~o�LP��k�΃��N~F�c��}��4�1���O_!�d���p��Qe�8#z��g�jJ���]�^��A�m��/��J./<R�Ǐʉə֪�jc$��bK��$+E�+��� �^;�FF����|���/]��A�dE�<��p.W�=�)�8َ�KKc��QQ�V��\�QPY�����GXl�t�Sz�<�8�-Sh́�J	������5�A�����eJ �ϣ����TT��E"�_-���,�M�H�Xg����t��)��l�C����>�у�_BY�]��.vb3%������m���S<��́�v�PQ�s	�`�����?f����u{>�t��95c��~��� ����ɉ:z7���b̅��R�W�I����q����؉U��+f�?@�A!���@dz`T���:0��9E�(��aF�+�'���m���4���r���>-�aΟ�s����;\�;��{v�?F�����PA��V�?�r�	�|7��׏�N�� �k2I1�f�F=�e��8k":�a]��V(�ڧ�n`��
 kB�9�ד�X	�h!���Yՠ�Ч'� 8#��Ҩ���X�ַp�me�����s�X��	�!K.��.k�����Q7��%&w��4[��`�(b+w�F���.G㾧mNmg����(82N�+��I���U����y�*X1�C�� ���[�)+�["��9�5�"`��-���Yx���2+�c�T��]H�:������@g%�+�bF̋�1�|K�0��=�M���y:\�4�;Na\����U������Nj}�n=lٳZ�;g��տ��	����U�/`d��p ��o �J�hט�sˍ[uG�o}}[���^��LI�)&1}8�d�'�h�����`�W�|��^<.a�N7��������\˹�X����j��b�%aR�y��Yhm���,�(���.�Nu�J��=C�^��Z�XF��śUj��7E����ֻ�=�l?%�a̸�O���*��	�Sz�Z��euZ�>�Pp�Pf�3ƛ��{���r��kI�l�cִ���mG��웯���~}�j��R<[8����hUY ����p%8<��S��/���,����v/>�+��]H���34^��YR�9y�L��c���J����拭'j�(��;6}'���eQ*46���4�CB�<�P͛�(i~��D�p�Ʈ�-�3V��ǜ�a������n��M�&��j<E ��ˆ̥;�	�}8��&L�o�a��r���9i�Kq��}A/������nY�nG�S1���C��>~��h�3��wۭ+�V��<�nw�^%V�O}r?�����=F}l���=c��<�v6o����6mq�~~iնg|�IY}P7�L���b�b����oL��' �{��7����i���h�e�񓍞��5V����u�;�X�4��r������{��lVn�h�a���7���9S����/�>վ�4].�u��Xd�x���1�֞�qo�Z;�k��2��=sN�ꅆ��D��yUa�3����|�cq2&���K��+�@j�?��{��+?��{}���?��^p���s)t9Vv[���Px�����*�Z�N*���\�M?-�|�=�\�%\�\!�v}�;*?���]�� >b&f��˨�|�uz�� %%XE�E+������
�����G"Hj��.��a������f��e�:�W ��޶�GHP�I�H7��~��G�ߌ��a��K�ú���UmkO.ɿ�[pl��o�h��*G��ȓ%L�
�΋K�(ӫ�^ˬ��t���j{��G�Ah�Ǖ��O>pS�3�E�&���v���� w��˓����Eeǖ�%�������J�*i���ϕM7OT1y�#]C�f�7������x���qo��.�N�g�O�<pf�Z�o��[��G�zOEJ�s��=�h2�%A� /�O�4树��8J,��=��?*��ed�M�X ��B�!u��0J�21���pF�����"
�[�}�Z��|��.���|�g��j���ۯ.�ݦ��������V'�n���J�F�V?4���o<9�hz��R��l8��ݞ�&�cw|�}�"t�^�}����UQ�;��ǰۅ�eG2����$*k^ߝ�׍t�1�I\��_���U��
_eWf;�x�Y�x�H��������]�18����S�u��B��Q����M�7�͚����a3o#JUPb��s7�8�����f�%�=lȎ=S����ns��ϛ��DV�YHk!��x�%�}��M�v�ͺp<?����F]8`����{�?P�����@ɄCk���ٜ��>E�C�wF��]s���� �>ʯ�D6�.�_��e��I��4\�k�o���sx���l�kG���^��s�hf����>�i�����Q��y��~	�|�F:g��X��t�Aߌ���-���3�!�]�zv�*K6q p�}<��(���NS=�,lD67���ϪR7|�&�=�hqxP����ԳO���҈"}�%�J�	�j��X���yle�/-ϻPJ�縷3԰ufƿ?ч�@��6���p��1�q��)��C�hno��D�I�o�>�}߅K���"��`z}��\�rgN�Ns~W�ckpOj����A��"�.(����ކ�O�q�Q���GFq��c���;G��\��a�A����-ԫ�;���r��;��]����b��x#���FP�8o��󶂺�6�jéq�Cٽ�_MBZ���ܡ�BW\Sj�9F.��~�`vq�
��c���Ԓń	�b�ꈲ`$���z)�^"آ_��;}���#���Hh�O������/������ґ�w�W����0�m\�KZ:��T	F�{?���ߺ������0�8���m�Fy�'O��i6�Y)�	NO��(�!�p��M��dt���EC8�P��7�;=p,v�����*�DK(1��uq����F/��U݋p�����X6.yj=����E����^���B�1A�3s짢��l#Jͅ&�M�M�z?6"�Qf�x���+�l���,Ϫڷ@ޣ�G	E��r��P3f����w�B�a��B�q])�	^P�H�#���r��~����U�(�Y���n�˘,I��<������:i3�{��m�HI�C�Տ��9	%�nn���}\�Q�s��%u���!E�p�u9�_������ѢA�^G�a^"Ȣ��L�t*G�cR=�Q����5�v'Sd|��LӀ�yx��a�8=	���R&`�q�)�������ٙq1C�f|�����\���L��A��a)3�og5q~p�q�s��l�l���!
`{S�O��10>[�Gh��bf�ݫ�� 1�!|�Ƴ�M�%��S��Eb�Z��[bC9�XG�n���oǨ� �W��?�g�t5X��ʯ��$*`�H��'�>
� c:88�B��� *93c&�۩G?����)/�����I�%�i���L�K��lڌ̔��ʟ��O�p%�ca+[���'}}�ZL��@��2��z|����Ou�����cK+/�T��c�Đ�Z}{6��+�gϜ�67�c~FР�d@�w@3���rQ��;ʟ�������IQ��g�ө��q�>�wPk^�?m-yw�?��bs.$6�5'k����N�d��P��K�Lf}���uw�2<oX��O���|��#&�p���|�<
 ���<��P%�Q�`�k8S*�27^b���g���,�ᩄc�&�Q�qɣ�f�����K���K��Hc'}��s3�q��h��
+8_�>��*�ٵ�ZWHphX�=Ｅ�wl=`�q�����I�J�)~�:~��;��M����gc���0��C;��t6	4�d�&)���웏�q鞻N�BgR��N�k7��4N������U��˻p�/Bj,'��N�-8u�S��X%5���Vy�(�p&=l�{�^�O�J�L�δ����[�~i����;�Ì��` N,��i#fzD�$\$�������ӝd�T��H0Y������0��d���9�8&� 1�!	�b�Z��t�-�4c0�hxl��4�����X�S�4����$(F���r8�o���	Z��^��d\�����d�N#����+'���l�ĝ�_X�]���Y���4h���m�og���x�@�J��]�(G$;��o�x�?���h+c�ң�i�(�����V����W�I���	�
��n��-�=7��ƕ 5y�</4gI��z-��|���]/�+�ᾴ�r�ґ�a�j�������*ڌ�g���=�=��1&(�w(S&0kq������L����O+�����݆	�^92DS�_̟�6o����� OPJ7�%�-�{��'O<�t�<2h�s�[�\��S8��^^�£��vE㲜Ǭ3����g2��{OG�����w'�Jg[#Ye��~�;��9߱�(bo�T>����������AteI�{��ٗ^_i��%(�l��������Aiܗ�^^~Zp�Z
�}���,k�jP٨�(x�p�|�O�]��� �0�׺���n.�<)ߘ�q��4{F�?p��FV��ڤ�V�/)�����<�bZE.1���ڇ�R�i]�����{m�0*/K#�H�%wRR��� �;�),2^hٴ��Ei�?���~i��e�V�A� �{:D�x�C�����e����vaY�z�`B��]�:�+v�.������C�1]R�2穜�|� �}��*6���z:,�����J h#��q˃"+�O�h��:u�����=����Nk��P�UV���N늙�k�Q�
�]��77ݏ�����0]Um*y��� �[]M�?��I�ܫ�����ڒ�7�?䛯DB�>���R���X$6d
��4������.F��]�erm��_*'��]��~,����	�ּ wtq�at����hll�������,�չ��ν���\���׉abU�伦G�z��v�Q�����}ǚ�J��Isz�h��ꏭ�[9}�u�S90'�A�6ָB���stD�bl�/��@��s�:W�Q��z!����,,�'1�x�Ս�rw5��9(Ì�\
�
Ľ���$��𽂡d��eD�ks��)��lZ��$hȞ2'�=~�[�CI��������pt���:2ޓ�4'�2����'1R�}£�-��B��{!X�����U�@3Q-"⍟_�/���^����U�63�c��:��jzZW��f�!<��}w�����F<��>5���2��p�p�l��4�n+���ʼ!��F�x�X]�sq�τ�9H��<ԣ������]&3N�H��(	c?��k'3Ծm��,*�9��
�5�'�D�A������WGaO��
�ʤ߯Y�h��I-*��E�f�"����2[�Zo�`�ma��|�n���[�xa��x�c-���Ա�ҿ;�Q_~�T��� 'j���X_'?�H����([:p�/t����-){�
�a�����[,�zR�0E�տ̱����zc ��9���n�<����*�g�1N�)?����#�!mi�f�]��$�>[϶[��t���Ov�Ȭ��Ɏ2�
}���&��cq:Wl���_F���kv ��ೊ��#���d�`ʌ�W����z�v��g<Us}��(X������W? ��v�wFFc�2��l���$��[�J񡻇1��"X�u����f�X�`�`�{�8�A�&I%��_։H�ΊZ���o6A�]��p��"ߧ���S��ў�y�F���о��Joe�Hj�G�"ǜ�r�0I����Ӫ�Ɯ�As��!M1��@>iS({��\����y�q ?����cC����-�Y�����ο�� �aTH�_`0P�t�!�*��vKi�yfD�	�ܙ���Ι�X��*H���(�X��aT?�R�(�֚��Ą�n��>֍�a�W��s��8x����{=��q.���/�s[�Bq�V)�
0�P��8����*�ƽő��:��Q�V��`2c�ª��Y7�#��x�2��nN������e�ڜ*5��N��8=����-�[�.����ځ�']��NgsK�'G~�֝5�+�e+�C���xx��ؽ��<g���_�8�����ꮧO!�_?�b���H��e:�c�amt��,/%��{�y�BΦ�������RǺ0�썥�C �� �8���N�m�W�	t�n��1҄��}�H�W���/'��2�X#H��Jl%$���$���M��� �u('&&�6�u����G9�}�<�D�$ϝG��ר����DA��߅�Ѳ���+>��S���-&�kI�j��9�p� ���h��M���L@}�����rԭ����l"�%��+?���2 �� ��� <���X��لa��-V(����	2�%�����DG�0�<���������fiH઎?�x"J[��XHz�õ6˯����m�t��c�P�`��ءdp���QU&�/�y$���7��Y��eu���B�_×#�?,���r���K��2@����j2��ҹ�Z/�XwB���YE_#�3l󸴻��A,���L�r���wC��e 4�h�$Z���g� ƪs]vf�����]4;�� �\]t0��J��:Xt�L�s�T�-�-Vi���[Di���{��Ƿ��(��Zc���W�5�'�KcV�cSD����|����K,��⿮ ��@�,���@J�j�TXpuN��>�
���uu�*�D�ú��XQ��qd�X>:����-�:�����LV?>&D�v�e-�#t����lH��eҨ�q����&{x*���T�,D�T�@���04��l�X~�F{�@�e��vz���t��׌�����M�+�7	�
ʑȳ֗�� ���(��-BܻA��R�o/e}�w�����C��b<�'O������667i�ũ��� w71^A�;qb+Ҷ�h6� z���J�����NAg(�He��������/A�br����W��a������$'hb�{2eU���+jߞ�q႔p���-�I_$0##�O�2��P<�T;��XC]�X:❕���������4#��b�_�ޱŲi��#�?�(-L�8o����%i iG��t�-8B����d�v�u��̝��H�w$m� �F"/!�G�G�o0#�w�4�j�:���y#�lK�qN�[2��}g�3�qȟ��5�R��U2�Vs_�GKk����DK�sz�ޒ�����U��أO@���b�b��M�Q��&z�A�bC\""b���6/�-�̢i8A����bN-���PF_���Ȇ�P��@F���"�g���Gm�]-	��04Sa���=�iLY��Ұ%���ҭ�7MN"��A
8B��Ӂy
}[��@vjɓQ[wyN��>>Sl��F=2x@�]sk����c�dM�'������N�����
�#�%Ħ��N�ܺ/ɏO�K���9=�!)a"H$��XL\T����q]�VQ���Z7�Q�;W��a�+���@\t�'������s��`�̾_�J�Nq��!��D�!@�L:9A��	����t�����0�v[U,����'U����.L��!ݥ|�<��=�p���������qd(7�I�H�!?�L�qd�i�/KR�e9��^/�Yuq�{�pŤ
q�}l;d-f��w�U|A,��n��a�?�O��3og]8s/�|ϲ������(�;2���n��xh�.V��S
���L�׾*��O������^h�m'�P%���TValW��Lj�a��(܈F�� 8bR�#�H�vȏU�&?=�|��E �&1���&�"@!�T�4�Q	�Qݤ���^~JS+��Wgu��A��8���5�ݶ�E���.Ӳ���!�_�m-��6�X%�M�u��R����%9>5��Ѓ��J=�ԛ��P��5���_G�B
_��G-�N^��Q�?+Dh�thk�rw�u���Q � Q���_D�`@������I=��dnjZ_�}�w�?bZy�v���>@��v�o�a�^��V�Ði�S�p[�3w�$��<�v��;���]��WD�e�4�����M�� ��L��E��(`��Y�)˱�Z=�w�� �����sm2ٌ�Y��?#��v�:�;D�7�h�YI�Z�vp� ҚW.�S7%l�]�vK}pA��j�8~p}p�vif��E��qpP�\�x@у�G@�W5L�B)NO�C�LP��NʓaR�����e�2�R�`鷤�=�MѾ�߮mEk���gn��A����+�B�OZ~t�)��5�����O�Ƙ<_�͍���}�n/��y����y�� "�%��"\�j�_#����ҝ�:�{7&�E������i��T��K�Ύ/đ :��w`ƌɁ��|�vT��*i	W��̸�x5�z3p��U�/�y�ő)�w��1���;��/z�-�| ������|s+����{��!�	�sЌ)�%�5"�'���!�Nn������Jd�ު������|���O�5�?ȮrLI��#T`�ǝ�B�$S@���o$.���"���>?��[�H6c����X�f�ۼ/�H�������3R{1�o'y�,~�u�PR��aR�5�M��X�&~��
5	V��5���k?~��������#?PWP� /x($�	Wl�X��tټ�'éx>�N|r!��7;"�w��F ;[/��g��S��&Nbjv�Cs�����Qf�d"K�6�cyr�	Q�P�0Ц��a����Ϣe3.�v�w	���:&���!ь�.��v#����&%��Q�W-s>Կ��	g�*��B�s,�t$%��Mߡe8�w�}���'W�B�)��\���$��>T�F��S8�]���T�	:�d�BO 	9%8�pB!((�����sfzRX(���g�vwx��r�]�'A�{���@�FG�|����u�~=���u��YPD��VW�LN4Ǆ2��~����ڊ����R�(�T`�V��(���6��֛'-�V�_�#i���$�Tt'&�wSC�g�P\�v��� �0vs� �Ao�3Rt��w��${-F��,Ʋ�ޝ�KQ������D�<u���|"FD�&���Ś���4炢ڌ}�A���=7���0��N/b�^�{J`Y��_��R�lj.	��
3��^`e7�-���ފ'E9�).!6�������pP�Qک��;}f�=Ďp�������}��92���5�.�
B)���-���d�A�3v�^��F4����)#�����J� �e�&���k���PeKu�p���-Gˈ�W �)�F�>e;}�|�fr15/��_#Ґ�`E!�U���C�[ZRAKX4�]��4֋�N�#�-E#��2>-h�)�P��G�e���yΟ}��� |B�� O�6�+�up�HW~ǔF�h�4���W�mSF�ϻ�s2��7��N=����F#;�Բjk�?uAw�J��u\�H�MW��x���#����j<oooee~l�TLz_k2��
��kX�GPկ�`�
��(u<�i�,�kEx��n2ڷ Vz���>�|H*!��\ɰ[DK8mXEs�E�g����zo�bX�3�`Ld��f�,�1�Y�&��B�b��qøx�jb�X<kgZ_Qh*���]���?���<�2mW��Z-t6�:[pL��z1�BDه�=������o�& @�a�*�m��W�;��!r��H����)��W���T��iU�=y,���W]~t���*F��+rj�e�J�^4��eH�JGQ�Rn�o
��W�V3[�e!�|�x��L��@Q�hhC,6(��^��$�.d��[t#�%�F�$&"�A'��s�֘�d��p�(�w��q=*݌F�{�N�SD�S�%͓����oa�CX���p���D�݀�jG�S�J'u�z]=�Iݽ#]}�:'�8�+|A��������G������d�)U�M�F��F~���AŕZk|8{�}y�߷��'���cq�I��'�<,	��T1��6��\�t�c�Q��,z�)4���,gKqB3��jaӐ�czC�8~��m�	��p��Eb���#"�Bϭa"�P=A��G,J,���;�H�P�O�,�<Pa�1Q멼?��(�c&�b$O��è07��Xi-n�.�"���,�;S�'�����ĕ��eW�$���Y"�-|��.ğE��XӸ�X/Ij�fʺ1P�CVƩ�5(���]~\��E�:��/�|+p��. �I���x���<����O3��x�!����[?Z�E�*�~����誷�ih���v'O���E"�=5V
�,�B�� ��T�)�Y��I#���o����¶��|q������ �!�y`�-z^�9tQ���$,DbM&�4ð��"<���7p�GT:�M�(E&�8�&��>�MA7?S�Z��E۹�T7>>�f��>������Al��-��;$�k E�?e�S��������M^<Y��X���Z2���L�_Am�S�XhҫI�r��.�9\n�����	��t��Km��n��58�ڗ��N.��o��Vל7�̎p~�W��xm���X��Z�6�x���;���Q$���*�,`�OLg�b�\�<�ؐ)Og�����7/F�޵�z��J� R+c}�&x(]B�`�t�/��ݤ����4��
�S���`�r!��+������t'����R.�Cѧott"e�B�%%7��,k�q����~3S�n�-��E�*T}5�[�6�|<h�F�(S��[�k��� *:��՛�55�S
a����W|��z�œ���X�p�8o6���e�ia�fQ�u/'O����:IC�"4�2��W,"�*�
?��d6��|y�@5�
^�&�I�E��i�ǚ�C�|Oc�PP��tI�nh�r!�gY�Viek�{�����R����"-I��)]�����D
G�b�|�l��4|4�����Hw�����%��?z���9Yg7��_�%diD9�Z�5��=�ލ�7g�j�[@	.5N�h���I�'b��=��S1W܎qԀ��G��*G�]����f��wq���ɿYz��5u�7�����P�ɞ9�#R\YC E�1Q�Ц�QXl�[��H�k���"�r{�5�#�nL�D�-m� K��X�1��L���v�]��X�s�Y�	�0J����|�#%s,؁�X���ݺ����T�xG��\%�^0�(��Y�c�I�ؚ~��2�Q��}�M5 �ٙ�T���ـ􁃉�n��~h̗o3�$0�VN��Mg�9�n�
�j���`a7�I�t�lY��}?�z[�|�c�;�L��z������rkoYi���\�����
1r��eQ*����sc��}=���*�R�=y�_�1�v�\��B-�#�=�R��u�1�\32�nR����\벻ڲ�����K�{�BOE(�Gd��լcC�.��:�>�-��DD	����/0�j�~iA�7[q}�HBd֢D�).*~����R�7��]sN�Mbϖ�o��x���xā�Պ�`���@ �5yR��=� �?�9`�2F��T,���9��j�I���d;{�Z����K@ZZZ)�ºoen.��t�������&�惱�1,X*g�V��7�C?j댔7]��2��E�	���
کK�G�L��5���{�Wel�-{l�ۏ�;����fix�	�(Xc�8�\������oͻ5��]x����2��ƍe�4�wgVKuK�w��z���*a���gd@e�VI������3��o��Y�ES�uC9�K�c���S��1U;!�`�Y���`'b�߇�f���?�����ǵ.?�@JKA���q[/;�O9���1N�x���k���ED��\����XzZ���B��n#�!݃![6S���G�E���F�<�eBr6�q$$�D����s+7ec��c��w�]3����.<Q/'���*�U�#ڙ�i(��@�v����n���Y{��S��D��b�y�z��*K��������N�*�akk�7r/.���l&�t����%�>r�a�/�,T������=9g�u���eq#��t���p"�~��{ZAC!��ۮ�:&����h����Ƿ˱5٪9L�<��P��Sa���R��HZ0�d��M���}�LȺ��<�=��l�뷖�a�����d�#*K���:I��qJɨ 
�l�,B"Z�~����"(U������E]x����iw��8�(p�fpe@,�8��X�Ą<������Ę����o�H{��o��$Pۧ�p�m�#�4"��
�鬙��\�AC��gd0:�a��!_s�~i��[�	�\����'��\�I�
	D�d� 	``�;�v�t�����9H���'�{����.^��"V.��B�s��d�i�?����2$�t�	d�	�|�d'Q�i��ii$�<00�adT�f��*�1쬸*>�S���j10P�L�#pAded�m��Q�Rf=��\u+���?�ŀ�M����q�%Gt�v��"#�"N43eB�@�Grw���k�����餩C�.�X���R�i��0�/X���M����J���~	�}�oaZ�wV��{�X>��1�������V]�������������_gdI'�C;͘p�@e�ՈR������ɑ,�m�;�����-[1,3�k�Nd ����䠐9悽x���nA&����f
lx��MfJ���E���3H�IH���f�@�^���|*�޷�q�:����w�
r56d(�+�������+�-�$��r�F���P���9�oU"��Ⱥ/Ɏ���s�ϔ���<?��z����Xj��ħ��#��&GN"�I�.h�'$�Đ)���U#�K!B5��Dd�r�ƪ�UW����=g� g�U#�r����o�5��] �oͧJ���z�7�1��n���Q�d���2�#���D�8ۻJa,�)����1+\F��M΄��Tዋ�>OVT�M\��@��5��H��`$�n��xPlC�T_"��E�d��m��*j!��B�Tb`�#�ʼ��5�"p:���է��b���@�n=�������@�OG��$�^���4 �N��x��Ʃ�ېY.��<����P�Z��S
�{^��`W�8�d2���L	�WN�#4��r!��Z��
��׋�b� V��y\!�0��D}��t2ϟ�J����[<"s��B��Ml�Ž��,8W�iE��H�E΁�L�v��]̼z
q�=9�`H�-#ca�@�_��Z 	`��3Цux~����t2I�S�`ӓ��3UϙD��E������OS������8
�\TX�/UA��<D�q�Շ<�����c�^<�\��,r�Ƒ���tR�qa[���q�ue�ߎ�k�}�'4|t����~��V�4q>��D�vJDz�X���T�ԊL@�"d����ORH�iP�����(�F��ä����el��hJ�i8�D�b}K����2��"�-��fD��diJ"٬Os��3�)�>�B�%�L�IsQ�ISG&��=�BL��Y�'�T�G��f~��+c�I�Se7	��B��y���C�j�g�
P�5����bk`����oE�����.7��m�lc�]�i|Q8����Mt�<��A8��`QI��&,l�ۢ��<m�\��uo��H����',��^����7Y���+�Ȳs56;;ћ��y��t.�65x/f�z8�`ɠ��띛I��=��Vj:m�����PN��⼡V��q Lsl��m9ZEq�B��1�)6*9�8�E�ػ`ʏ5�Y�����du\̓�@V�6<�ްD8�9�dV9����ۂ訨�h^P�=�� b�C�?Ĩ
��D�䟎��<T�q��J�׋�og-�l�Yv{�����m��O�
���T����K�c4�M�UuvH��F�ϼn�����9��\N2��Xp��ܻ�r�B�2����otN��7Z"s��||��FF�1��OW ��DQb�=FJwe54�Q���t_��@�$Ĵ���H	zɽ��:$����-��W\n���=ye��Iߑ'�F���kZ�]�Y�1�8QH2%�4� VO� �RVꛇ W,
�]M����>������r�"��rs��j$| ��bC�����<�r4tb"��I�0�X�r�a.l��4�9�~���>Zկm=��q��7+{���Dp����rw�����ZIe$��cs�����x�d�	�3��L�)��D�0�]~Ƒl��i5#��X"-�(8�ߗ�5��!�UP( ���X�Q ����yvU�(4�UL-ȉ)U]x��j`���3���P�y�b\d���
�w*"W���6Ƴ둬��EM]x_�Ҟm��D��e&�׭��r�`���x&���so8�^��ąPi� ��m�G��"�mϷ�jc>}�1�ntr�#�,1��1�\'��檏��4.�x��mnk��8��A3���4�orw��̉k{[�C)�0���� �P���7=��3�\�)T�z��P~�A�r�3Դ%|<Q'�`N��U����R!��s ���.�Aى?�E���m i�Pǅ�t�B��I��9B����X�nc�A�41�7\�9��%��\��@�Y^� �aA"H�ǿ�*|���Nbfw�sm�7*Iii���.�Z�ֈnC��j6Ⱥ�;~|A�n��>Ξ��k ��:�x��p��e�bOZ�s��OZ���&h��J��Z� ��B�0�q�<�2����8铖gs�8�K�b�%�"-�"�o�ٓ��HFBX?W6�7���!R�@�VX��ƈ��H5!�?E����2�]��+��� 
v��M��MWUUmo��-%�ݍ��Hwǥ��^@:E�� �ݥ��U�.�����7ޏ�����g����Z�6	�����@��}kn��.@��$	g��� w�������)���T1jf8���z<��}��$_��p����'#�20���q���1.�J���Z�C��.��/=����䠾3���oᄛ�z����?C�1�O���y�vG�Z���T���E���N
�Q�D	��S`��zq�)*��h��#!�X�h�-��E�$�6fz촔q�����)-.o9_��3�T��<��QT!����ǥ܀���r�4�1�*O�-� 
Я!�z_Ɋ��M�`�h|T6D�HT/�,CoF�W�ۢ�۰�X$}L5Js�@�#n��7oF���1����� �Y�Mz�|�
�Y�(�<���yw@�����?�s���`S{ʳ��ڰ_���M�Z�d�XJ��X���Y�Mq��_�I��
�b�i�WYԯ���ig3L��l^��#>�A�O�7�y]7�7���̞ɳ������IѼ��+�� ��x;V��B*��?Mk/0�^
)۵����ƨ���/��� >� ���v _�H��nSB+UA�;��P#Q�/7��!48rmmd�h��I����"G>��m?���Oi��`�3���tB�;��ٚF���Yٕ�39����K��8xpr�H��d��LK��-��p9�N��xj5|)�±�����[8�7څ�BE�2��q+j��Sm)�Iq�S3�,8~��ڄu��r%|�̴�O�Jϲ��Z�!�af !к_�'��3|��߬L�=� lT�����ji������3��4�۞���X��Ks��{���/.~u���^Y�"K<?�����O�s��LW�D5}�ȏ\��,�^�@t*t>���0)68)�R���\���&���1���ir�}-����nR_�߼�f�!}l��I5���Ú�]+�����{B|eSUK�yn8�V��a�@��8�ޘr���"��ֶ�C1)!E1�^$�����&PG�KE��W��~o���h?GVe�w��H^�*��z\o��<x=��8e������7KzYJ�
����&_=:���S�'�^�
G���+P�l
L��~:��Nw�����h����l@Tgʃ����:�`|c6B�U�yz^ʑp�N�23�1^;_1�';Dh��	�*1|{keD٤����P��rjj���0�ξ��.�/;Gȭ�|����3�6~K�K��'�h�&5�z�ә����E��v
ml��ڬ�Xw���}pD���q�g箙"^o�{^�V���ڃ��f+z�į���d/=3ju����@L�K'v�������?�6���JDK��)�}r|
�Ub�y��כ�ʜ�͋�?%�I%f&DO�b9�I��������l�O�aT��t����S/���A�ۄ�������_ �J���D���]��ο���<�W��5��M�Y�o:V�Z*���.̻�����KT>tq�F�A'?D�j�8[yF�q��	FaWe��r�z��/�����m��I
��J��4Ρ����-���]IW���tJ�
.=ݻI)��g��H��!<W��c�?--������sma���炕E�n��2��p�V����{��U���HI%���&	ؔg��e�s�Kw �]���w�\)���s(��*Ώw[����+"s�
1�r�U�mӑ�0uEw���[����U�����>�$�5�<l>-ːXx�ur2���,�\wZ��^�)uAYL�\G���U�e�
fE�n�~������<��I��x���bѿ 9������0�I�����M����؃��R��|L�6XY$p?}� ���k�«����)߉�˪��Q_��Q��_�7mJ����q(p��X�ȐUO3��6\X��9s�?��N-]8FԵ!N˜�����,8?��W�����QĎ�����V�+jeYZ��<���,�T��X�>!��U?��Ǳg��!�$���"(��B��L]�!����ƲD���* �s(���_�i,r>4$6+����Q.���j�Y?�x�˳���w�q,gO?G�a�u��q��N/��"ft5�.;�/IC/���&D�h�/���F�R����,�T��m;y?Pi��ܺvr}���,������C�-K���
�'�A7� U6Ӡ���%�!�i��c_H��uuYEM|���_��h��A�&����%��ęF�4���k�0�fa�1��˔������wA���s��A�wf�$[�@��
9 �:�X��d�J�P��� _��>O!�
0�6��~�"��=�(�]�p@��Yfs��Q� 	�e��kwV�#'��X?�e�A˕I����L�%����3I�!��M����@�9k���TaL���k���Ի"l��r��$޻=&E�W�GȞoG��!�=:KG��gJ�D������6Ԗ�M��{��jE�WzZlO�׈b���f].Q3��.���Z/ٓ��XZ��g������ޚ�N7�	_+���^n�}8�"h�}Z���'�\��eЂQ`�h���nf�D�:�K�0�*��Y��	{k��,�;h�^�E{C�|p��{D�p��y!o���ͤ��-u��7
O�Q��j��Z�4��ށ�J]p`����͐6���H�k�@#�B%f�g��<a��_�7���f��Fbd(?t���o����Ǡ�މ����Du�P���1r4�G��� �,�0��0���'�\9)�!�YP�� d
�fI��4(У3Ã��g���Ҩ27!�����0܍��[Q���_>��� ��Z`_��m*^:v^��?��\UkL�0.p麚�����pԼQq�����R~���tB��z����'�8��]$AN����Ͳ�� �锹����IO"w*�cQ�I���/��}C��/[�7���쿯TV����	M� �?�v6Hq6���?&ⶸ?]AD�x6�ME���t�;�����✻p3o��}Ť����rw�0��$�$9��|řj�.�?����\_t*��8�[1t��t�9�Yˡ�P2S��d�v5c��}�R�h'��yҬZO�o��9(��r%R��,ſ(��13?���"�8q�g�Ds�0K=��`SL�qL�GG�.�i��'.)L��X��8�'=�r�f�Bf�ӑ�޼�O
�k&���_ɨ{"��X�ilQ,FM=g"k�t����@M�x���Y-��P��'�OS�9io$L��1: -[�k=)��R�|aȜ��H�}T�Ag���b�:)7��Ϛ���6� =����� ����vfΚ����"J<�.��-�x�r��E��v9�gfrj�i�d�1�5bz�Լ�'*��Qr�Y�m�H��%2�{�ѫ}C��,���#�Ͻps)}2.�ׁ��!�>VL����f��1��\p/���o-1&� 7���ǽn���l�L��d�,��k�_-��f�9=�	�@Bɼ7	���3@z��n�Q>&1�L/Va�/���c���#tk���YG���l�gc�h�NY"|��u�bKD�T�1��m��ꊍRq����� �t��p���T�����S!����iơ�A����t��K�M
��5
����>�wQ8^���\ꗍT\�p�P�L�a��c��ݦ��P*���t>>���E ǴA]V�����)��|ؐQr���U�����D9oHs�d?�i �o� o~T�O��=������+^��cG���W�Y�J��KARH� ��| ^(�i��R�IW��y�I�2���՗g� f=�(�g�'g+�k���S�x��!������mO׋.�Cu�괉�]),�q�֠���0|`�`�٢K�@��-^+�p���K�z�&u>|ja��aBcs�ǭy�D���6��?p*,������֝Xu����1�ь�;����S誠�I�&hxQ�m�z�j��$��Wp5�#c��;�&���&���ѹ&2���0�0l�� BLԋ�	�2��!J���L1��uC��g,X�7�F��^��W��Sqۛv}V�j2�嶘!0;v4Ӳ�R��B�#ìk��N�&v��I{+�"��p,&��&��Z�Q\���"_��M%�Xz[��?@ylӪo�
{/j����T�>���x]/��c���mjJ�A�~���G>�p��"�m�4mA>�(���,*�`K	"8.���Y�$�g�t�Ƴd�8�"\�<�ݦ77��t?�%^��-6N9ڱ�mOjc��1�vz�A�x*�x�V퇃Q�EY6},��x�{�zu���7�F���o��ti�����*Q~�`�G���a'ZL/Q���$���g�������zGpow-׌�����*%�r����+"�!��A�?����L��ȏ7)�~X�;)ؠ$�0s�1��D9t��-,73$^�q�0�!��[�PTG	��DC���i��q5�{T���ٛ}yP�	�U�#s5�?�� ��!��&O�[;#
}n�
幗|�	1n�u�8&�Dv���Ά&ڂ�{
O�`T� �ʴ�?�Eaym�����7 �E���ю���87;�$��,��"�cZvv
Nwa���-7$A����߈R�i!<����ĉ�?P�5�.pr�JV(o�����)ܹA1��#K̮Q��x��*&O1i���2��s%�W�<�m�ǳ�-��mҿ�ͬ13˗}V����v��v�D��*)��}��3�[����D���2y����.є�W���d/C��g&B��q9�ù������!ޘ�Z����X��Ʌ��]��?%���,����wi�rx�c��Z�Mt\����5��[@N��Z�^��s/����1�8K�I���g�~�T���&t��/�j������۸Q�T���^�e�6S��Z�F�bh��A�xx,G�(So`��:]H�ny���Є����$�A�>Y�g��2.���̥>��v�:�K��֫ޏ:������:�KX�@��b�%5�Y��DQ�����Z� ��rՄ�g-�E��:N^�]�\,G�K*�JFe���p7�����?��N��6��j"{��-^ͣ���oS-�Dn�T�[��J^|�3;�x�[E��j�<(*UF�A9�R�~���س�����hq���w8�:����*e�,\h�6���*��ed�f�ڟ�Mj�h���~���r#Ml��Oִ�J�����!�0�U��bx��ۋ�'�(��v��IĒ$�����Y#�ÛlsO+�A��ݤ���B���G��O�V��
�`f����Iy������1{t���>������-�&��Ǹ�"�V��.���_fWK�J��
���>*�M̀(B�j�u��vz��R�l]��3��.�Ls��c��d>?����zg+n��S���ű`k/����3�v6H�m$=p鈋��ĥ"�{v�gyH#���[�r�m}v#�&Hg7$��f�D����}}�JnʜW�?��<*'�bee��#�M������\u$A�ɥ6]�rؐ�O:/b4>�Q>��a�I��C �q���-��Q,g2��΋sz��T�����6��늄^�=p���F��=ʻ�'��!��L�}<ۿDv�n� � �>��i=��/�c����u��'=>�f���#>�q1'��ǇB0�.\Ƃ�\GQ��O �H��'"���
T�Z 
��C�?WH䛃����X�t5�6��cv?p��n+��㈠�5e*���c�r Q�=1t�R�\8ɘb�|�9���?��'d���i�� *��;�h����G����HM�./�l� U�rVv��c�iS2K�)+<���������9����"yھ�jۨ���LhNnS<ہ�.��Ο�񴧓t�1���t���C"!=��n�aE�Xd���K�?׍�!'��C�t�dIc�#�t����ˑ`��ЌF4R.�����b��0F-̺U:������H��s\x�ܝ�z珶0P�T$��q�n���+�f�Ƚ.����^�w�V���H�F@*.�"��}�#�����ؿ0��`�f�-��kc}UT��.{�s����xE�n'"���5�)9���<=�g.�u-�6�'aiu�m�/u��.��XȢ�?O���lqo��Z��em@H��g�!�銟��Is���1N����Or�(���@�ެ}�������4��$��u�t9Iv��!8���|��X�������%�4M���C@��Tn�П������P�Y�����`��շay��J�>�Or�����a�p6|2nb9��a.?`X|��9��,)�vp���9�t����?T�=Σ���� �\�����̏v���S�>���1,1��p�B+k�LN�R'2m�E)ѕZ�-Vw�p�^�5�ZV�jJ��\��%�|���y� �ϧ�����|�8�=��O�7�b��`�@t�ej{8*�}�~F:�'K>hԃ���Up�1�X�!2�"���L�ڋ�����=���q���n@$&��SI	���q��$ѝ[�k�;0C~!�tӢ�<a�4�b�_��}JpI�j7�� �210䗛���zo���tE�Vj7O���NT�x.Y�@J����9/O�y��n�%KV��Ŭo�L�C_�\a!)�����w��rѾ&?����ܑr^�h=�^N0�ޚ��j��Ls�#ٌ#�E�(�؇�?���q��??K@j�s������%2KWI��$��خ_�~���|ר�.��3��^�{�6�E������=I�N��P���97Y�,��}ة,����� ���6��`�����O��)-�hn]���PT�ю�\�t����u����Y��o�6!���[�n�vqH6��&��-"�Dq���7�!�V���5X$���
CX�f�_H6e`� 	Wh�&�X� �x6�͡����
g[Yd�L�� ݍh^d5A}��
SEJ�L�!c�'�P���%a5ZI��� �	ޛ��aEK5!TA׀`���DJ�V���F���q�SZ�M�9�H�+0����Eb@����-&ğX���דu���pN�O��<x]����f\��xX�A��a�{;F��f?Z=
.ue�T}$����W8�c���Z<4��i�﯉�G�L��>�b�h��$�[�����/<�D[ۑ���L�2�t3�g�'�绝�����}�u@��܄&��=O���G���)�;a�����>_\tc�Z����S��t3�+(����1��40d{|����R���I������d��`�H;�s$l�/0�M��gL)��E]�I��ς�R�rX`��������"��{{��6h��rT�J�jg���؝�6���u_�Hc��$�b�D�VkͶmGyL�ZP_x�*�\(0���	�}I���	��$=�=�{��� ]��M�m+��z��v�B9A���.��-OS�x!|��^<2��q�`��v�v��V�TJ+�Ɣ��3���:��U�穫����L�P/��.��;`������M����қ��{%�t5�*�m&Ӝ�θ���5m���h_�_��W��Ofk�U�A=��y���#�M| �EZ}�*��Df���{
^$�]*qZ0*�1`�
��	�ݞ� ^p����!��V�X��~�,JuA\��Bø�l��eTƦIc8��",͈#�a�����orx�s�-����f���8�R�W1+���I.��ͦ����Mw�mL��׮��8_0��\X��(zSO�)��f���u��|_kb'���:���z��V 뾘���36ӯ��@��v!m��g(���[��]���*���X��9�_�匉� ���`C�6�k���R�D��F�ҥ-)_�|��,�F-�_Ji.��3�B�p�eo�j_�SW	?LM�;�Ejy�]y�ȑ�k�7�58Y��; ϫ�~�,�rx�0�c�D�@�x�����{6(�1'��^-�G$.n�����l73�W��!����L�1V����~�u*����g�!1 IE����?��;��8*�)R��,I(m<�| Us�N�BR���NLf���m�IL.|a6-n��%Ɣ�?bx-C�btԝ�>��b���~�Ƚ���8�ŠI�CmA���dR�F��.XY���\���z���Q8z�$��]��0�H�N7~�p�����3ʰ2�ܚaXZ
����f��K�B�Uf���E�,Ě]�[ l� ')�r���� ��?����ә �<��F=�� GmƟ�X.CR��(�K87�[F:�y�얛��[�o�o�J������=w��<l�2$�p�7�_�j�l����N�DE���if�w?x�}�`�a����Z����������dM�|��8�J���� �d8���б��)��6L"�@��g	l�cj�$���>̍-�rs��3�GnR�-G��ށhr1����{*Ӆvޭ]����z_ ��
h�>��o��U�-�8��q�*����}����s�w:ha�6��W��Ʈ|�Պ�X��cE�����Ó%�'��#��C�TJH�
<��@���d�u�b�g��5��ޗ�U�'��<0d':m �	�����Y7D�#���D$�?o�xv�������TN���B���#���K�d��-�!ܐ���4˗oZ�d~�C��GƁgJ}�0�T\�R�IV�K$Ӵ{yv�����ќ@GKKK��x����lHH>H3����.9$�����7W���G�0�㹢�X��Q�?��&$
y����@��m�����1�A,"�]@!��K�)�+$��/��R�O6Iҝ�orbt�,�o��öAQ��G�(�HG���tN?�~Z�>TUd8۸�P-�����Ô�KP���~���V��2	`��9�m>| r{f�;���`O>J�k ��f����}c���}}��N�h�g^&�=L즱�F��J�8�,E��N�����/�y�E��������>,��Ӆ<���(�vQ'�
I�>���3�y�ƣ|}�%z�����{i�?�2�MTH���ɳ�=��5^��A�B/�pdTIT�:	����'�`�7�)I@�%8m?H�c)ϡ�J�%3�"Cw�T��)����]����!\V@�����~���"�O���T�Iз�YL�C�����-"�/
*"N�0��2֒Ԉ͒�6մ�b���cX�3��y�8�+�.S4@� Iڔ<u2��&Y�l���3wC	�.���Ȩ%�sE�Zt��G[R�����NK�1t�٩_�d�C�����,p�/+,{�PU��� ɻ o�(Ze��_���徢X��v�V'�:%4�����m����t���~�,��
���8+'*��Q#�,}2�x�E��N�v^;|�ͥ"��o��y�[c�=�����h�{��ƭWB�dC����q�l��}�	V��\I%]�-�@O���R�D��o�Y8#1�~�e�Of{�5��A2[����'/��U�����c=$��A�&�����R=��x&/�cøͤ�1VV�t�O���,���g���O_��Ɏe�2��w����+p�~r�4L�Ι�m� 㘊G'���5{S�?�8w��@��"��7Hԝ$F`����Q������B1wI�lR��7<`,/`�������D?�!7��ܾ\[p:<��#�m�ř�}q_�ӝ�T��-���+
��n$��O�[����Ҫ�Q�/ߖY����ҟ�(�z�}�AٍXQ�����h��D�c�����½�	XY?G��!
��d��e�O�#���9p 9�T
7p�S/��� ����E�f['����rp��_�@s�y:������W@�xE��&�TB��!�{8���O�!=�Ff��૴��D�˟�鬘F�߶�႗�~3G���e���\�	���	��p��T<NS�_R[��a`�ہT)b�}��p~[B�L0�cJ?"�|����Wg�ӻ��55)u�W� p��S�R�6h4Nr���]��v��l�7���MB�;N�%
�l��ٙH{���e���m	��z�=u6���^�O6/G��
�P \���܅q�"r��P��Lt�$c7�OE��	g_����ٛV����YN����̅[GV֢�a�轩��R�q��Q*�Z/������늗+�f�|�F%����x�us�J)̓s�:���@ķtc����@.������C�ވ��,�m&��ċQ��*��M���6!}��v�K�U�4�e�U�#E�/Ԯӝ���	*���L���5��ȹ9Hi/�?E�%�|¨����u�xC��mvS��
���Vu��S
�K�c�n�`�>�m}�2��6d��qPc�����(|���5տW�t�8�՘���n��=^:���A[��jE
�3;op\w]h�����϶��ڼ�)���Ѱ�X��1Bc�\�}$]��M�zߥ�j����Ė[Q��n�A"(G��v�j�O,�������=��S_�.�	Q��D�b7o�~�>4���]�,?V߫�UE�������u���?B�ۧ��}�������|�a�4p?��������Px��M0�σ��0[�.�#��XX}
���K�"i�����ϳ�m;8���ò��]�A��<Oۢ�ш���N�@^�[����Z�r�]�Z�ۉ֭kY��h�| ��Ӓi� \�D�zV���QDԚ�&;^���g���i���.|��}3�X(�;q��Py��0�Z�f�e�ϻ+D1�l�W[ dP����|��5{���4'�p9��T���ǈ�5Ex��<9�3(��]q �nl_���j�[�]�/p	��&���|\ʜK���fU��������?�9f�A��s.������9�^�m;��#T�D\:�P���������C�x��J.�:Qt4OJ<Ly�nq�IU�������Lt��T�f{Of�]�-雨�>��T>�<+���]J}��������p�� �Z��x�r�U��M�'کr�:�����:�`��ua<-��
�=d�������/���ڋ+�5d7Eߋ�K;����$ KQSMTR�*���@|�	q|X�*�9� �CF�4�����_�xw�S��:��b}v2��X�G*�Dj_F�sU�B��~����h�&v�i�KP�:z�@��w�r���0��Ѕ&晿�'I0��"|ĺf�����II��'j(oz����2r�+`��t���'�2����s��U�!P��6�Q�'�x���4�#1����}R�\��F��.�ȯ��KF��t���I�ԡ1	�#�̑0(�:	g!Q�ޕ{�2������!_�p$�,�f�w���5��qR�����!�mҕ�j�xx�Jݹ�U2�SY|Hb�A��0�Cq�6/{��x���;�8=,z���/�_%�?!���gR"��I�N�I"*��}�Zr��y�Dxp�,-�R\�8d��|�C�7�&M�ϸ�oO		���dų*MT��k�k_-aq���s����QT�KIy�^>L-�<��x\/~c�����S�ƞ�o}�V8O+P&�g̨�`WD���5MAr�(�4fYXR|m�]�Q鍰j�_ �����#x�����ĸ{�0{L�%G�����Q3���*�@VVR�������\�3mgD�����p����ُMϼ��4e���%��.�.lI
z�n�v�����z@n��|�8.�<k��N� q^��\u�J��t�y�yѻ2���(z>X:se;�5|�hg��	��C���o�*f�Ug�r��-�xZ�c2��T�=���],�aݓyv�/=��:��=�#��%��ɳ���;�R��f�\�R8��G�y��������*@�+��m#J
��1M16���`X���/|^/?;Èn���k�!؋��i o���v��/u`"8z�ˉ�}�*�O���D��%�٘���f�S�Ϸ�k������z�[ds�L�P��-�����l�R�1a������~/c�!��r��T��Y�ޏ4�mV7�0k"��M���%���.Z�`Pg����H-<�V�--:�� ,�����pm,�p}����^$	9��sEo�4^�$J)�]�Q�LG.�B�簱��Y@����I ��`�T�Y߂�Z�h��Bveb�,�ha�q9\�.��m�$ҹ���l���}�~��b����a������u�6i㖖�%����P����h����F廐�X�IRՙ��Oa�}��X��q��hM�ϼn�Wy�q�I5�|���o�v")T�rO��j��uT�
��R����B�JSz��!�v�HF��Lڳ�=�N&?��<�[Do�Ų�I�����v��H"Ä�qlz�zz��M���o��Z#z��.��M��i塢�l���T��1b�/t�<	/LD�-�48E�O���Q�4������=Ę�<2)B�#%8Ky�MM�:2�Uyùî�d��m����yG�L]y�a��#��k�w	��CT>Fu�N�c�6���M�u�$��[�j.����U7�'zum���5�9X}g�~�S;�C�:=7���4�/3�G���%>@�W=��<�Qms��Nؑ&Q3���.)���?����,��Ozڏ_쳓|ڠE����D�������X"r��,��J�t?bY0�������X/�0�p���Xz��v�~q�$Y�r\kp�C���vaNF���˃���P7�i�>�~O���[K���F�_�g?A}��$P̭̩���M?��m�7=0K��B��;�ߐ��4��g�}|��4���k#eRއb_���)���M��=���"�꣐vYJژ���N$�Ʋ�d��%I��#�<�'T�����e�č���/V�z�h玐� 1z�צ~��YE��O&���	Z�y����U����Dq���~Ϡ�j~/�ӖQmg���OoѸ�b��bi��G8�S) �)�7�#"���_c���iQ��Kj�Z��i-$��@];�6%/�����/hz�d�],�&U�[e-��R���*`�ʶ}��AS$ߺc�<�S63���'�6�%��Q����ږ�T0u�ݷS�rF�I�Q_�IqTR~<��־r!��B��_O��C�`�L~�t�H	�ϭ��he���o�������nq���Z;hq��'����6��w�2��x��O]Baj�"�Te��=O
�P��U�o��T}f�1hz{��(+58�+G8�Xܧ�NLQ��.`иN/�07�z�LشP7�+��,���f�P\i�ѩ�jf]`D_��ڏ��ׇ�	�W����_#�ɛK���G�,�?8Qzg��^/F,΅��/ܔW4BH1�MJ	Fx�έ���&�}�w�f��(��Q%s۔����'&��O>:�m/�F�8�5�l������t��6����J?L�l�ʇA��Ż��E	>�g烈�:�%iZn|�r�+�[����@9��Hbi�x�[�Ͱ�{e�נ�Nǻ^��1/�JoD�A��׻W�ЃcԈ�����]����o�L6�H���))�D�P�x�mg�MX��%9�(�t�K�J�JYL�;��e ��� P�1f��mǄv��2/l�����G�H��&]k��j}�s��k䭦t`W�o�{ld�YP�$�d��������C ɹ�z�Z��6�iQ�|�=JT_O[1ʹ�5�9��h����U�"��	dX"��'L͚�yF��CR�(,�����J�a��$G�UN?p\��y�U�jOK��`4	���Z��. \T�d늇�|�(iIy.��ͤ� �&��@qK�<��+�����Y��}.A9��a5�:� �TMh!��%T��WP:4���)�=�:B�]��UX�GD�Y|4�7�;&@�����k0��&��]H�e����H:�V-y����9����B�5SI����5�,<굸\~�w5�g5��h�� 50G;�{f���1��~Et��{|�	��$�k����G��r�6��x���R�vgȆ�~? ; )	(֣��){tB�zp�9�-���~X��a����hˮ�����gzZV_k��	�]���J�۾O]pS��
D�����fTN{S;DZ����G���{������,~��>���qn����rS�'�F.@�P�H��psinr]��Ʊ������g�s����xތ�5]w���.����l�t�3��{"M���6.UǊ��}���4��2�.�2��fE���p:�UxT|=��?cbE#���������\�P�J�k-��,6��%\
�w�f��Y�Klё*�����D�c<��uꋐ�~�[�׺Ƴ����g��i�Q��_``n�C�8ra����w��'�sM��lP��l���J�ׯ��~�����y�K�)b��wݓ�m�#@e@�!xs��#挌��7:���]��:��턂om��.?w�R>�fc�>c>y���\�vt�-�LhUW-We��?�ý�����-
��<q�Ӭ��r�����i&k~Y�a���bx�� y���Ә?4��9D~R���]��`��w��	F#���D�Ǳ�Ѿ�9���0������`2J%_(�@�5|B��_!�w楟6��(�b����sʧ�?j��/^
���p�M�L_w��։48�^�HJ����`����kuۗ(��Or(�wC׵��3�ak$�QX���ʠx��o
�q�I�Y�B.KO����	�v���z�v��r]�9᳥�jXO�l���߱�m d%=t�C�������y������a}��G�iau�N����'��eV�ߏ ��
�z.{�߆Q����u�o�6j?�c
�� �E@��n
���Hs���,+hA�{��u�^A�Wm@x���7��2�lnV��(��cf���vNcJwñ0<���%x8G�����q���#+�Z�:K�sː|1#z��"���M���p�^3����ë�'?�>Tx���i�o|�nn"��螭:�o��c�LF�����k���cc�3��a�w������j��*��e���6���z�����M����q�!4��gNlפ�4��.4!����)g���k�����"(��_�zƺӥ1���5'�~x�,�PT�j��⣥8����9,�,Y�p?d�V�̤/�-D&`\���p�46��M�U� sڑn�����T��J+~m�U��fp��툼x���0*!�.~-�"��X�9�Ae!���oA��M�ܔ��sf��WnV숵�D&��w
eX���9 �"(��@�7�*K�e$$����k�!���½�/9�9�\<��"�"��0�!�磌TU/q�\��s���ndB.L���uQ#��I��q̓Xr��rx���C�U�j嬦�m
�����VB%��@��J���AC�=[�CKj����V!�w�,�������4d�Li5so���5���,\��/�KE�;)������㽳�&$=ݹe[)�$@����DG	�k,�����՝r��tr��^�>ayڮ�Q��e>�jl]�'�M�5��
g��E��'Iɀ����b�CaK�B�N�3�l�����S��<��k�WU�\&U&�'�+����Q�ҝ�?�8��E^Ko�!�zV����m��"�[v��v6+$oN�D�mQ��-I���ߡ�P�뮜��̾tPQ�� ��q�0�2�{�@����:�"@���I�`�j7Ku �|��4�օ#dl#�/��p�}��;�g�����<Bd��Q�i�Yy)�E�&#��S�@ȼc�\0�Xgȣ�#��n�39~�Z�顇9��N��2(T�zp���q�����׷$���3&ŵI�W�[�.�P�b�OO;z^�+�L7�-� cZިJ�&V���tHc��������Ƙ:�d�5�s�Ǧ�W��7[IR�� �8a�9f�����3�x��ɔ([�[kr�&_H���,��t�����S���?�s3��H�z ����^OK��N��5ɶb�3%<�IR�H�{j��i�ʚ�����~2	���)��+��<�jz��`�������x^#wa������^��'���;��/�+6W�C�s��~��U�>i	R�]�j�lhy�P�dSt�S�'>Ρ��+�_���?�񾭬�qYq�j�ϊ�H�����55���[�Q@���_}FѾ�8B���*o�%��1��m<�fخ�)�Y���]6��R�qA*u|9G¦�]��{L݀��,���U�����t�"bB܅%gK}��̕#].��㧚x���񝨀 �EV!Z����!�*�ں� �tw7�t3��42��04ҡ��5ҝR� !RC�t���H�����=�����>{�^{��sf��?lg5dr��˾�EUm���W�5�3���L>@�~���c��Z�&�	D���ů���`֘��&��=8F��&���)��p�3�&�~B"��}D׻��� ��yٚ�Op�ԟ����b9j�x��(F獫VkW�3a���tj�:��o��mUz���x�<!+_}�������&����B���w�FU �����*��
�:>��O1��ʱU��>�#��w�:���y���Bo4H�d��x++r�%$̶�Z�Ϧ���_�\���W����}��*���y��������&p����Xzk_��n����,�i�5���hL�Lx�^[��ƀS���C+���ayl\���*x^�E��Ʃ~FG@)�}FH�T'���|�ݲ����{��u ��ĺ��'@�N�[u��WpztaL�si�A`9\�)�%�(k<���貯S�5CW�Q��9��JN�V��z��T��q�5�a-��r𙄠��h Yh���O���9�!�G�@AlP&�H���f93��8}}�
�d?,h����U�7E��o|\��������mL�Śac��"!���-�����  ��Lh�n�3��|�f�yk����=�	�hq�����J�\2 �b��{�ɮ##.9c.�]�%���Ⴀ+7b!�HE��&5��r�o��5�,ş�U���r�W�ܪO�?�^���F��� =T&�8�4�7��%�6��}���zFX�dz� �U7$6�f�g�G�36hr���I�H�iȗ��������y��>�W���?{�ߙX��dۨ�pU� 7���s6�-��<�z#��e�/���M��W;��8��+��Pk��B"��w��l��E��"�3DD�{�� 41+n�(4��Ic0�b)�a��;J�i  �z�N��zźI,>ߣvd}��pVY�Œ�X��}8Q��6���	��~���t�'�'��0�9甑xe�;z��EʀO��T�,v���Ӡ ��"���>M;ނ��jU��yZ��b��w��{��\��������E�5�5�͜���#s��q�����f���vV=|/`;����r2��Ie	u�b��[{X�caK������0bg#���s8�������Z������ 6N�N*	��cL	�Tfͽ:�,�����	�Є��θ,T8��i6�[O_���1߳	@6<�}Bצ�T�N��˽�$���­۟<d�};T����
��4�W����'��h�Կ���/�Ӑ��X��%j��,��(����kx�i�\�`e�`�eC��c[cS�mg��K2�I��[�G�ōi���ꇳ�%��4%�RHgn��N]RXl� a�xQ��!��\쉞,�m(Q8�Ż/m�0bl���Y!y�������O��r���@��S�,|\
�?��pB�]s$-��K�j|�8��t+��.1
���i��&s�zW�p�`��o{쭵��#�����o 5t���u�&@܅ƾ�z� �C	����1;g���2At����xڹ(ib؀��$h���LVXT���I�I�ʔ��"��-Z�D�%{�K�u���D2V�,����>f0��'�t�(���D�Q�Dv��5��~��7=��f%W�)joW�ј�M�3
j�
u�P���F-Sm�?W��&�!7՟'i!8tt.;nd����bL�������҆��U���&Y�7��wti+J��?��As�|,��碈�١�}��C#y�Fj�[D�SJc������Q��a"�G�����j�wYa�R�t��=E�RC&#�S,1�Q0�zh"�-=�e�(a��jJ���� ����CQ��-�9�����Sw�e�^(�t�gUr�0! Є{�)��"��U��Ku�i����%�N�� F��-i�O���޾�$�����7�þ�A�7�eV+&_^��DJJ>�c�Kc�i!B8uE~� ��r��/Ъ���y�Y�'���kM���?�����}F�=9�~Ȼ��8�^�U��2��������B���Tk�q��Lꔐ�����%KM 7����l�ܭ�V�N+w��w�abՌ���2����w�����޽�AI��t�m��Y!��H�0xX��g��
�=ķ�j�S����	I���r���8�-�c$yWp#I��N�12>���Yp�$��[�~����]���/���;4���ii{Z!Q6v'8�`�Nve2��d��*).�y�S1���s�C<o���pA��!�G5��0����.4���wb������9�p������޲���+]4>Jz���Ӊ��eX���tuY��x?�1�!���rh��4���P��)x&k���"�x%�Kz6���/��'|�C�[[u��M�^V=��N�r���_R��>���62�7<�_�ך�v��t^~�����إ��np�]C� �����I�������u��UF��㞿��7|��m��5i;�s6H�� #��k��\���kkJSK��Z������n�$�4���/�K�nJ�7*�MvwiT���}º�3�mZ�j@Mo��:\����'�z-Mq5�����A�o�eq9@�[����"���)X5H������h�#_}�f��Kv�kB��zI*m=�Q	{Z�l�[�^��<˒�g���52���A�,1:wgu�|]���h@r:Z����5湷��S�/��a�l�y��|O���"�F����&wt盘�D�ƀ��zoy�x~>��D+$)�7��2�u$D6�� ��/�i;�"���q���̘�R�k���#LA;|�y���_��-�p��V ��4�ƹ�デ�@�J�fL$^{��/�
mO�7V%e^�d���1�S	�N�%�F��S����4O�TQ�n�?n|/y��d����tT�5���q��ǻ_Ƹ6�'��_�sn�,fIl�dj��hu.O���7�?�h�b�C�T�j�lqK&x�0VJ��D��_BF*yI���$$P\tYJ�n^=9~��L�T�+�2b0M�Hbt�|�m3����O!m�^&�z���*�]��b��n�c���:���U[��V�`2ͅT�v{�`�`�C�a����bx�ֽ���dk��s�!l��XB�v%Z4�P\b�U��|*��I�7��1����U�{G�)0Ԑ�9�E�+DS�+��jS��_%������{X���osy�<"�<�[�����HԠ&�V8�����z��.|�5�L,�#�D:0��4��Қ�^�qµ��@½F>�D��<�S�=>��)}�}#˕�L���L��1�:J��~9{YaH瀑���֙��Dؙ�=���E��uc��; �ʖqS�媺6���Bf���Uw�X ����;��J��XL��T�8kD7i���p���܉�Ͼa�w)�ǹI�^���佬��\�5��3���.�3Z��"ޠ�d�M�"�_�
�Ē��41"VLj�Y��>6�+}*����A���%F$=a�slZ���L�=L�zq��'��'���Ǔ+�X� ����1s�,���W	F�2sr{s�\ak�c�ꑭ�*�gF�,����F�rg�X�z���v<�6C2y߿�>k�hw&��Y~Z6Tk@��������Mc�/��-��}�28��A��UR���"�腃�Px�������Ӛ3C��䇅��!!�����:I�:�����!ʾz틅��-������:X�H��^Hz����X_׵��P��#IQ���o4�&T��+�m�����&ѢZ�t`��ƫ2}t[�o�&��=�N�e�E�X��V����i7�4���;��e㤫`u��s�I�k�C�׈����#��EN��!q%��}D����S�����RκȤS���UC���W�4�C�[JK��Y�;V�GHN|#������� Y�Λղ$�Ec���m����1��l/	%9Bm�7������tSA������lH�'2�6���dp=S�rA��?���!K�����Y���Ӊ̞�__Lz��~|(����GfY�ؗ$t���V� ̅FG|��~�V�xٺcy�s����w/�0..��~a�+���b��5�:o�M0z[0:�01e�IvS�m���=�p��c_i�����`�/�g��r���<7I>%�wG�����ŋ#��U֌�6�oM����4մ�9��TL��19ж���Z�_�L�����͌v�� �VAէs��L�Z��d�eX��"c�H��B3�������qF͋�������*f$���͔�cֻ��}���	q�q��n�+g%�Tx'[3�t�7w�oH���MU��g!�Wqlެ�PS��*u�U��Ͻ�u/�%�l�\��wX��	1�xZGo��`/'-�x(��]q���&"{����7?+SJ2��Z\:]
���By����/�Q�
�����{�Z�d��v�v,S��'��F�fdt�3"�#"[�S�Yw������J"w�>��~:�c-��?+��J0��3nNϘ�Ҫ�J��/���<�T�f���ܶ]1�o����e�ᲁyƴj���D6Pi%���Y��x��]F3٧�-�*�T�pWNH?<�%���8x����Y\ɜ'���nC�g@���i��� [)��͎���yEt����/A[����(V��*֊L}�j��n�+W2����sf�������s�̑�3 K+r 8���-~Gr�(ukLӇ2�F��r�'��w��'B������vn��T���������]���M����B���7�.~N��>\���h��ڿG)Ǫgϧ�		��_�y����g�ڠmm
9���7�PzcL`McfKޅ����~�P� j,��~B��ev�^>���'K�_�˾i$v~���0֭�%��Om���o�E�6�K'm�������*�5]�ٹ���ys*�5:�.Nm�OLlտ��5�n�Q$�#FheMD�G1��&�t�T�&�qs�/�7wp�]���S�v�	3i/|>�Rz��"�l��~��$m�N���Q,�72n��dUE��{G�������W'O���;��͖Q5�,Vf���?ގm�k�l�/0�zg݀H�m���y�&H+�z�}�&1�ƇO����b+�b~[�bw�eVN�Tg��%I1OK&Y3zհ�����zm ��d+�����gBí�<I��}l?����f^����G�˱��G��q��O_$�M����6K�Cmyl�
sw��78	/6>g�4��'>��`�Y�2�"ʭǩ�_����T͢��	a� L<8��J-�z8]��bC�ڤ�L�;�8��0��
k�9}��C��������z_��.ʛ�y�oW�~��ep��.�pyB �y��?�,J��S��2�ڃ�M�����}��E 2d�䫇�ͣC����6b/'��|�m�&���خ�+��&.�*哧��l��}�����- ����X�w��|}������۶�>��j��b��~��1<�+	e *�8f��1Mq��g�<"0��yX��ֿ�2�)Z&��R"AO|u��\�km�n���\`#NY?���7������L���������r��V�.A$N����u�w":C���M�b���Gv�72���6{A�a2��U5Páw:?�_Ӆkb�r$�͵��`-T@7ό�V=���*�/p\��M���WE!�fD~�Z��]=}菇��R��&;�29�����1$E #"��j�xY�B�aG4i��$��-�М�6b��c�V�#aB��,,�|��r��49,����jG	l�`���4�O�ql7~�6s��v��u��a�u���<�P:Ā�z�_���v; �K�\�ؙ\h���u����]��jO�[[j'ґ�ḀE7F�������ɍx��>m}�p�|�U�H�L���0����S���ڧX�;қY[:si
����r�sz���_{T����sJ6�!?�iȆ�l&��U힪{�)u	^=��v#U��`'�	�tUaD1Y��=�;���3���x#g�s�"�&�$���وsjp"��f�	H*�.8W_���A*��Þ�N�I+;�)���xN4�֌~�>1�O<'��������v+K|A��,g�+�3��Q��4d&Ѿ-.���t�8�pё_�Ҟے!��3�)��zY!�>*�{�'�_������@������X�c��Hk�i�yL��v�#g��.����_
�)(�?��Q��L���Ax��g��c�c��$�b��s!�N��+B��>^
���Z�����r��ɺL��Oxn�K�9嗒�{?M�Rs�0��w�tD/���3�d�-Om�q=�x��sh��@+/��0��'�˓z�� W1�]�D�c���d�;�k�	LpL�`�ۚ���L<Z���-��ث�!�&�PG\��2<b|v1"F���~���5�h���/��J�y�S"p��Ӹ0�d���Ҋ��{C��B��9?��@uY��z%�vm3Yp���"Zk{��������H+%W+<���b��'h� pl���������'�76֞?1b�t;�LM�*�Ш7����Z�X�MͭjŞ^��5����'�]ْI�#Vdp:Y��e�{O�ݮ졃ƭ�F�~�z�\I��vQG� %�3�"!"�ښ�V:��J��A5�U(9C`y�i�����=;$BY�)H8��y�I�L�f*�U���_�d�Fz1T��YB���!�/�u�Ҵ��5M��Xc|+l�~6U`w�*�2�җ��̝ǭ��p��%���|�CB؈�쏗���j��O���;���?.:"��7��ȍf��i�{By:��ү�%g�6��M}&K�����/=2�J�;���X�	gy+/�L����3h"�$$`K>��L�dX07�h��}��`������1,��+HyHJ()��ۇĦ( ���|dZrh(�t F�&@��,�45�-��H�1ڛU���adl�k���d^���۲O�+d�MKK�"�U�/�U�ꘜ�4�����ܪ�-a�V��)!��h� ����E��+�'P�/1��`�ZnJb�X���R���L�k&��4�,�F���.&�`���=�^x�4�p�5�� Z''��'1��+�bٓ�T�XҢt�1����ax���_1@�A4
�j}�^�.S���a�4RD�C�F@aj��y8����Nқ<�T��ΰ��Є)��vBh�2γ��<��EM�R}���Ԧ	eu	��Ϯ�w�u�(�0%'��j'�PER*�Ȫ�q��93�%��l�)�,�~��Ǒ�Ub���NnقMe=ޮ������$��9Fw����a�sI���`�s�
>�������ޚ�e���w��:�@�2;\�J'�H�|i{�hNX�1� -��v�_�-����}���	_ex;���QYZ4�� � j�Է��qa��*oGXTF�T(��c9g�-+5��џ��5T"���Ц��f��+�p'�6�ղ���^����j����]=|�#M�u�5wt�c���b��Q,4���t\�
� i�����)6h+[������	�� ":�7 \���f�d�[���A��k!A����
�p��gu��T�7�jǸV�o��ہ�QmäZw+�pnTm��gnOT�����N��5g��$x>�5¦�W��ң8ƚh�PT�#8;-3��#\���T�P#A��R��H��Y����L\/ʘ�E3�Bi���F�����3�8����I�j�ùl���0�,�z�(z
�A<�Na(���*Tl:��ڰ�A'AaX�s��ĠRǾ��v�1S~�&�]��/;���l����j���9YmO�.u`A�IK��I+����x��2F�Wэ�!y]���O6����b_;r4��.*|f ,Wz$I��<�)��h�/�3G�($��&��:@ٹ�j��ڀ߽8�y��e7�����Su܅��ҎHH�ʔ��ӵ���ܴ�4Oc�S�Q{�'N}�!Ϯ��IY��Q�(�5�U6��A�ꆷnZ�U���>�ar ����pR���8j^,��L�����c��f�b�
{��CMr��0k5h�(5Տ懇��|&q�'�l�9en�vO��+P�n���;�?����79�г,mH� ��	U��"�|H��M�S+�J�|�ٯX�7�����r��z!yem�`��V�/�iWi��@�`C����&�2���K*��c�r���q��^������+1�=�?�����{B�/PV�2MVii�S�:��<,U���h�GeԐl	8��D"D�Sa;YV�H��X!��P����|7�z�m.;[V^7(.����^��]��2КYT�t_�t�v�8�D�ը��KK��	A���r�\���#􄇏�cl�� �`r�zZ�pJ��@򕰭l��zI��Ls���P����.�_��[���@޿�P���n���"j�ì��ۢ��K���y�/�]q=�gN(d���[Q?^}&�1�wE̏�'�_�w�����s�~o|�0���m=�B����n�z#��I�,#��,N|�g�	lYԚ<��j��Mʰp���S]�i�f�
Ӈk˚u�!����6�U��҃�G'�a��F��Y���X�p�o�@�'�U�ȧN�9.��L�Ƅ�$:��
ػZ�s��ױ���I�)xtH�����Z��>�sV��솮x��^��;�4.\(���K�E�4��eƬ�qQ�Ѣ��ߓJ!d��TV�lı�Q�O�ȑ��6�ٛ	�0�}Vۑ������a��geV�bϱQ�[���':���[(+�F����^9ʜ�f�*T����%����頓�����CI?x�5*�U�)fB�%_5beW�}�b�+��3�~�(]����/���Y!���XL�����n�c�Z����'�3j�
"������'��wC5`SDG ���=������kW�	W`��,L�o����щ�Fr�n��������rN�����Eb���?�N��÷�kT����]��m�o�ѳ¢ʐ;��\ݥ�m�`�V���!�]��.şT� RG3M���.�U�Ө";�Z�e��*��� N���K�?�a��CӐ�f���U���	� �g[T�*���'�	��AB1 �N	k������ �[~Z�R�j�5�g�%66�M����Wb��cK�1���1�T�"WC�1������oq�H)5F�x{�o���$�~������h���g|Օ�?����j��z���'�6�4�}�{��э�"����wo����ݹ�_!�b�,�d +�п&��c��h�˟b���k��K�O�B49�E�lJ&���R��Z\����6h������c�	qqk��!sM���(�1�w jy�?=We��5�y���{p���y�u�����Ǩ �RLe�e,DF�&0�Y��>P��J�3f�`f9�$V�+V����Ї,̔�B���R��\���L_�'M#O�J�a����x�rE�!ӱh��Գ�?}Ä�b=n\�P:?櫴�-��ۗ��u�'����량�-ǋ�[0��Ie+���E�� ���]Wp���I�a� VX��*��x]$��Y��0�R�Y��k%�1�/g���$I��E\5Sc64}λ���(�C�bf 3+rYxmI�J-��������1�ԟ�⛢�Ӻȧ�j���d�3����OI���žA��^�>{���T�d5D֒�o?L��t6ȟ<�gu�a�3C���7h�PsN���ae3�2A<���N�#�5��&y`�2�wd������j �$� �z/��m�5��!D�:���;�H�w�8�S\U��BVE���&h�Q3T���e�W�� c� J6R�UDJ1�]�V&=X���Z�8����Wb4���¨��C�Z!����)Ք&޼�0���	��������u�(��8��>��=1����)�I/��!�� �V+���-�D�T+6h����#��X��&�:��	� ��pR)u���r �� ��~#f��o���76 t���ǟ���U��(�?7�a���H��J�gLmH�pPɿ��؟u��* �pQ5,?���Z������3R�V���A��WM�?!a�E���x��+Bh�J�E��9��d�%�Rg��c�<����ѧ���cԬ�̢���'�Y�6�r��d�o�q(��$J�)��H���m���no���d�$�/�Խl�y�t&Eg���r�+��I��y�ii�ժ���Á��ckkk1���_�"����g8ͽn2����np9���ȻZX�4�xo���x�r#�cֈ{��v=$�������/rމ�4����Z�$Z�c�2���2��Y ����,���禈�Q�*�T;/�O�wJi:����E�~n���qPzF�� n���9}�DFj�'ŏ��{q�;�vڢ�"�t�Z�̟��ˇ}-#�K�į��K0V���t����9pcE�s��;�ÆkQƆjό��Yc��M���mN���*������6�*�d��j�xd�@4KD����#�;r�w�<��!���Z��L�8��W�ᬪrv�R*9J�/=4s,���@RbN����� Ȃ d�{�|����݌IC56����� Dy�)���o����<��+lW�����p߾�(�"��6F�`�WMɿS3�	®g�A�0W}���}�}d�p>�x|_U�>~�۷��"b|�3V�ؠ2V���l�۱/����|�8�$Bp&pmUQ"_Fu_<��,�Z�1�[�^ ����SU����q	v:�����VB���nF�yb� ��ǇB)R������0���2���V��@�n��E��?3G�6�-a�M��փʹl��ȴ�t�ԏ3o�?�6ss�	���p�����T���M���Kh������:�����PCF+�F�Eۣ�q��8U��v)�:d����1-i�0�V�0��9l�?������2���D��q�B׃�\�F���?�{�:�
ce5i�g�֔��K�G��a���[�Ԏ�XEU~e���Q�:ae4U��O�v��o|�[;M�#P�F�^ɨ��6�e�`3� ӎ�h�ums�E����-�3���}�O����㇘{[n���ٶk�ʻJ�8Gk�0fvE��(�L!E�KF�{&0�&�H�J��ް���Ea�����%��^�k$�6�28�!���3��kv��T!&ǿ`�� �pD���O6����ߖ����~tF����X1j����j�a�Zr�q�\��W�Mb~�����2O8�ߺ��㋧��q޻< 0PRJ*�\)�^xPm�����Bx��n������*��XY̆���%�08V��ZXe��uV�|�x���k�.I��Niyύ�R
�I�ș1��Z����<d��X�ֽ8�c��,�*�O+ {��{�h�@����7c똤H #�QD�M�u񿼊�%!��ca��-��&R>�>���\�,Q�V��2�$�5�Q�9�������������}�06p�c}�08i`
�")
���B�f���~}1|p��w0[c����?�J
�b�?����9��g���T�P"�wS�3�[1?�+7Ѧe�����C{f��Y�I����r�+�[�������f0{�(+D��ڐv�F���K�P��@�����οy�Bmݙ��Fԁ�ZV�9s�RǓ���iQ&P��T���a5Li��-U�'w�8v��������W�P寪�R�o�w\q�8e���u�~^s��q k�E1�T�|��7T�RQI�Z�=a�x;}ݖ�7�QdS5��_a��XE�pq�B��'�`�6+Ģ2B�/x)�'���cd���C,NՍͭ׹�e��ڛ������G��K��+���*��(#�4��y�k 5��S���l�&�1a����6<�ia>ht�EӅ��o�sCmRӬ�lj�]'� d�
6�<g_�o�!�Th/LmL�좋�������>Й�������0�⃎�A�ŞH��,"ąp����l42�8-�c|�m�Ԛ����n=��\�]ʕ��̮ �a���\�8Ĝ6�A�S6L�3�]'�k����n�
�����~�.��~{ہ�ŝ2��3(�{��w�byy,���IOM��;�a��%�LlW��i�Q�q3U����f�l}N������x���*渿�O)y�X1g�w�o[9B�x�?�p�?�A��(���J3��̍/y�"*�7�6�����e������=�:S>�����r��>2 7Y"��}ل7���dS�L�^��5'5���`����Gk�d,̴D�b��*�	�����|�ϔ�������<�ƛ�j�\���NKG'�6����<�eڈ��5(;�e��r[�y��R���ڇ{<���:�����y��?mR���ps��
��䕭���.X��ڤ���÷VI�8z�(7)˔a�0"��F�q�߈���H�J�3a�_���"�T]�J�+o��{?�U�q
ȉ
�U�v��e꽮,�}\f �a.�T5t�؀$>��?k�_����	(36J�P|��,�mV-���|�:��d<0��T��U�w5X
p��j"�&�5�.z�������I��0��J�8�$Rɥ���j<<�̣�$8���!I��ΰ�>saw�]��� �T�����}�\l��%��B�]����U�0;~������;[_`�P�mGF?�g'Փ�����������t�Cm��}g��O��%�>i�1�'����N�����d�zp��(��~��L���/��vY]�ʅ�`���Ѭ����uKr.;~5�?z�s���oz�d|��}�#r?��FijX4�\i�!��"zO}/�p��	�!Fu����G3�:s<$("M�VY{���<��@�H@gtS���ᰩ��� &�#�%� i��|>+��/�D0�Q��3����u�Fi �i��i�ЗX��_x='8�s�z�D��!���`��vٔk�QT��6�7P�{F�"ݚ�l�N5~�v-~dl6�N��؏��m�x�8I�<	m�,s|�s�%�v�hz�3H71C"�Wʟ��Yf,g�{�~"A#���Jx�`3! ��Bmhf��ӽ3�`�'ڸy8!-���7�-�'��S��O3Al'�� ���7���;��f�?$���Pk=���=���0d���n��f��wz�{/	����T��Nj]�P�0���������X�3o��k?�'Q�C���#�bc.>��R"�I}}
��4���=�yT���e��d�{1��?b����6���b�x1�n6j��X-E,�"b+-kƓ�z-��˲�Z����x��@�Q�[�\Z簫�I|��8�u�l�1�3TL	��x�`�c�T��x��N��2�}����@*��t*;Ԡĥv�% V�W1r��n�y���@���󷋷Z]�;D��+&�}���m�w��r��ә�{Rׅ�M<�;�F�SDDj<lZH�`��UU4�+>�??y(�������^�W����I��o;{C�llU^sNǏ���X;�ځ�ʸ�����'xcH�Ygu�*���>�o�D ��8�������|��#]�J���=�%Zܟ��ކ��'UxUk>v����	�~�bû~|s������J����sl��YI���<�:��[�j�X9T��۷�-@�n2J�\�mck�����h1���e����0t�W5WJ�����N�I=�tU^B���!�� ����(�W?X��T�����D.��}!�)0IP���=/�z�ߖ���[������+sr1��l���4�������7�@�_�R�Ƞ� ��{%��X��͋xd]�����4��+�5�Q���IC/c�?1Ϟ�9u��,>�A�B�փ�`��V�6!�^z{3�fB�o^89�>ħ��_���*�x$�$���d>C�Z�����M����M��L/�5-�����~��j��~�;���P'[u����P�`�'����7I�#y����/	��s�ZI�z.����j�^<��i�	�/�L�����������~��Ү6 ��p��%*�=wOHN�!��z�@g~*�A��Y w&E�`$���w��C;[uJ��:V���0�V�+�,3E�?��aX��g̸S�/!II)���/����"��W�X�iY	�_�����$�}�
|�ǡ���gK:��nEl�(4i���H��
�YqCKlT/�%��L��q�Y>��(�4��4@G/r�wX��#=?NMP��٣���v���r8K*�"=�\.��WR���5��,��"
0"�ǒ��pn&W���<Tz-��STT4�p�b#���4��C��V��(௓k�-�UI�q9~��F���._��%7�4��e�X��X�\���g�8�=���̿e�@�Zm4{�Su�焌!Ʒ��)�Dq7N���ژ���<e_ȕ4+u�M$��P
]��)e �	������H(�w��>���cc�ۀܤ���8/>��^_��)��B��|�IQ}T�g)�!�0�i�e���+���/\�cQ�\�mJ^v�ξq�d�:r�ʮ� �Dxr�&+d�o����)m�A��L�e�e��K���5�e�@0����UU�ճ���O��lᅺ�F1�8+�O��d^���kَ�&.�e���b�,��ժ3|@OO�!4˾S��%�!I���*�V)�A���o����.`7#!S�Y.E�O���s����	+��&���2��b/�(rD]-�A�D1�T�v�<�Q;��Ζ�~Okix�~n:���k���e�R�@��&�9D}�U1$o��|h PE:`o�y��t'�P�0[�^ (#?�e�ڿ��5�j��K��p�J&��Gz"���D�C�1��
�T�_��m�a���g�/訓<V���a�K����v����V�#�O6ğ�?M�4�/ώ��*�լp]>��	�<P	��=�x��`aФ*�H^��`f���Y������R� ���Ь��=�"BP���J��0q��V2$P�����@P��ULO����⧈����ڥL`��J�K��r��� �U��2i�Va�c��#�s�w��6m�����o�'6�~�ŝNq�D�O%��N$�#]<�n����o5�t8cu���=�$�+ �&��?�|X��}��9�Wx�?��n?7�{��U[��l�W�RGKc�~~�U�B�3/Pe�� n9\un��t��f���P�Sdo_zd��h�@����6L��%Ԓ�[�$�x�	�������3��j���$&-7D��ⓦN��}�Fdޠ���aA�`go
�y��������S.�d܄o���1<��vbv7�ct��|��b����l��h\��L]�IZH��1����SP��jf`3/���I���h�BDM�߽�����@N~Z��Uo��3��sP�]cc�\�>������n|�F��а����2��ƽ�Q!��W��CE�������j[}nA��gŊ�b>���~�V��u��ۭ�ֽ�1�+��\��O�YSu5��x\��;�ĩ	�I�W�n:��z��2�
ċNu|-��~1�y�l๎��:�N�B6լ9.7$퉸�y�����`" ���Y�W[��_����e���{��@2��?��\�|X��fad�%���n���	p�siTX�An��qX(M*3 �Ei��pO��	�?2:Q�˿���8����'y��Z�w0��j�k���XP ��u&�8�s�!�*�R�g����̶4FT,.ź�gv�~5`�k�A��N(�?K��|����$nsz7Ք�!�A'����4z�Q��mcՙgK_�8��yG�1�%S�4���ܒI��������{�ߩ1x#��1�o:�^�,~x9��h�H� �~�gY�q�BwNd/_�-���Rw�*���~F�z|�Y�м>��&��ic��nsz���a���*���&��֐`%E�u��3��<�$a���>sZC�i�v�A�� �DX�,8���D�0w2}�P�1{;�����-ad<�5� �p�w��U���I�㞊�S"`� ��v��.�i�^����*��� FG�A��;R�up��r��e�1'Kv�&��ic�mdH�X�4�o��s���;�^��,#�TL��X kl��` Ό��,0�`�c���
Ì�rD��]�/M�P�^5��!j6�S��\h�`^���͍��O[��0��'���\iPF� ���9C9U�d�6���6����¨c�j�c�N��J�b��)U;
1������SX�(�r~7A_���	�4=�{��.���0�ȫ�]�a�1�A]�d�O�d�*�q�:j�'/0����t�R����f
�&�߲�K��{�i���)���aqO�� �CE��lX��~��1'ʌp����������y0�K$��/v�͈J���Ӛ�p��������/O��������W.M���b#]��6��!�9���,������)���*������k�����ŝ���H�w���Z<w���S�x��P(�@�;A�Cq{���{�9_�=[�Y뙽�L����I,0�b��Zރ�������Ƣ9fl~k�D���;,�,ر� ��#$�j]S�.�_���?���И����qv
ސQy�����	xs'u�s��ҡ(Yǰ|Q.W�ʇ��z��{� ��$�zP��bL�?�Y�=��N����*ؾ��OI��C"<f��S�$/��}@՚�����C��9ܬ�~�ceI�%{�"��kDůg������:���
����\;w���GXд�	Ud�%��5Q��gH����,��ڥ���,:�ͳ +��Y�[������$ipG�^�w�D
::!��
Onr�!��`����%�԰,�J�0ݬ,���Ҕq�X�֯��/���3�Y�4|eű��i<4��S��699��4��%��߿��j.%E��t��5��$�mn��~�Y|��aɏA�W���U'��G�Ad�{�U��a�������a;��쫽WV��Ǧ��s~����Y�!�<�k�V�*�q,,ôs�?臣ȯ4Ѕw�B�jF����ku�2�p��:����'��[9� A�ros�ݯ>���-��T��׏CI�;����$@S��rmB#���`03h���ow	f� g�X�pH5Z������"i$�H��ݯ�آ�Н1 ���J���85!+���s�eVf�*|��EZ� �E�ў��ӜT@�賏a�T:��e� ���F��5��tf�GF,؀��]_/I;L1��h��k\�+̻ʏ�;�ä�t��qm�յ��T��Ċv�/
?w��a���yULlWd��[p(h6v��j��l|<0Z:�~2~��������e(���3Ɨ��괘�S�ē4����Y��Y��|Q\\�t�|��y��6/�VAi#:�}G^�h	K̾X��3i=��Q_����7*�Խ��u&�v���pK�U��f�4p�mʪ�:_�D|[��#�&6.uV6�����1C���д�ly������n���g�eգ�����]\�� �5V;.g)\N:��x\<p�Q�*ˢ��^��Q�1i���g�CWo�I����d��>�B]������hEd��py��=]w;GÒ�,
3��"�Ķ�w.jk7�'�l�	7BG�g���[�����,�|d��n�m>���u?.u;�n����
�	`�o��<�7,)�yz*S�ٕ�G-� ��N�Ǻ�_I��J\Pv�ɿ�h{8[�/���%�y��(�w������ffiˆś���?�D���2�cndu�a��8�[�S,���=�>�!6����Zj���5E1��=n\��g*��b��-��O�1�Y��OhӓOo�r8:���O0�_��n�nN��s���'z�	���~�;�_	��\�!k���$F[�)C <�-OIH���Q��t=bq�E$.%�+����_�S����|?mX^C�C2Y���nDp���m�WP3�(-���7¯P����x�yB����-�*i���.q%$&7g��[����������n�U�T��D�c����8V�}囥�G#〳��_A�c�hG���"<��w�)����f��}����:0�O�Q��(p�v�;�1�QQi	�4V)�-�=yU�v-�Lm��]k��d��ز�xh��;�Aw�����VDR��d\�-�����7O�zx��H�'Q�������c�����G�Νw���н��*�|�cD�7��tk�'�'%g�am�+e�(5 ������ɳ�������a�`�&W�}G���j�M�ZB|��E�s�]��UK�c�����Y`�țt���X�Z��.χ�zݱ�����8�nU��5�t����0��6b]-��i�Q��q�&3Z�2��Au��(	%I���_uȅ^�_K�$����y�,x��q>���X�w�-IK��䃯��z"����ѮW��|$�3n���v��HҞ�2/d�������fse֊V&0������Ë0�]�Z��l���a8^89&H�c�(�JG{�U���A�@���D��Z&�wx��:!���|�l��?�=��Ԭ�q����.����e3K����B��.���q��Fm�}�������{�v�b ]G�ϭ쬢N*��w�Z�^d��\���2p����`��S���5<�(���S�LlO*�����y�b��]��*-�/�.[�^app(g�A����nf���۲��e���79�B�u54����gԑ=�\NۙE����+��GO�ׂ��9��J�Tg��T�v_}*|�l�B��d���5a��}�T�Ӹ
����fD�g����s����^__�M��]��ի[��?l�6�ਈTm��MT0H�7B�	!y�6�����k���v�\�l��j_�~~<�8���)=<�=^��q6���e�K��70���.�q��y�% ��Y۩e�~5X���f�j���e=+�ġ9���m]�R�`5�?m���n�<b�^�����q&���~���{�RL&��0�,e���T�����[%T�����jY�ʸ�LyS�v!U�k]���!��^M�L��5'}@&X /���^������,ތ���@w�XZ&�K�'l����Kx�u��b� ���J�5"(�4���G���*���:8���dP$� ���w��O.mu�ǿz�ނ�2�Rz�9���E�1�_�Ѣs�r̄Q�'6d� ��{�q��mͿw�%!b
z����L=�=��28��7l�:�D��	�3�6a�c��C�u�:y7ҝ-���c���.��V`t���.�F�+|7�o ۤ�Ad���*ǔq�+�ػ�d?n{Eق�J���H�0xd�Q�SA�X��A4���Q8��D�m��@~����a�94�v�E�y~ގ;oVhV�
I��<vǓ�<�l�5.\S-�<,�~ۊ���}0��Xt�őe��y����j���٭0�7�S�$�=���/Q�a����"D-a2,�@�I�W$��% s~�?cCLnzF��X�X};�'(�mg��|\{]i���#�1�䨩6�f���٠�|>��fPL⪾�R�Ϟ�j�U�^gT|bK�¨�q2�-L��6\�?�����q�2t�ܚ��g���x^�?��ӝ�.��}��B2�	�i�0Y��)6���)�t��eA�?����h��%~����v���wO���L����|P�� )*Y��u��Ƈ�b8E5'��b���'3�ešv)��E�6���QKi�	��F{
M�pa�6b�ynvN���gxk�T튇>l@K)�d���o��>�����T�=|زKFMf_�(�������(� T�W�|�8+�ٱY����\�)c%����e��1�0����8�bRrm�`�U���)�����_�l����M{���
�_/���� ��;��̉�ߖp����6��L����)�u|g�< 
�L>�w?�_Y�៤b�ng�%�r��� +��^�^J��>ӤzY�����Q��m������ɧ���}��xxَ�`�c����[�p>,�%�͕�S=*�xr�oF��)u�4�Ha*��I�,ۓJ!�h�TU���b��ջ��n#D�P�QC����y�j��l5�J������ň��.�[\����e۵��6K�e�����Ã���U�n�K�C)L,���iql��,��ά�˅;�%9l<��=�q;jV�;�VNl�(gN���	����_NeU��,Y65���CY�F�r]b���Lm�ѩ��B�����l:��"����P?�-��O�Cߠf�8�M�
�R�)I�0)NL�,��O����3����s��i�n��r�t��A۝j�}��۾���%�#��:~����.F��z��m%X��4n�٤s��T�G��y$��ALh�V[�ߞf�!?8T�]z��,v���d\.:^�s�/J[�>��}:������Zr��Aq����
g�;��֧@�����xy��O=�L=���(��x�ǁ=��\K|t'��.���au��8GD����C�W����=�}Ww�c�u�sy���î&=\��D� ���ÄV�m��0~Y�O�a
ޟ&G^:��9i�2�Xv� S=�kJb�՝;#Ңj����"�erAa�.���a}���u�5L	5�AuPf��{����Ogt�S�����9���?�Ă>���-���2(���A�7�˾��;�1@M�=�����6��O�Bԏ4�@4O+]��%��Ρ�/���B��%����C�G��*�7�6�ϋ���>7�ll"đ����Z/O�۠��d�����t����~LB�4v0y;!Sa��0&��C���qf���ܳT��V���~�α�_��w�׷�__�UTK�J�xw�/u]=K��)w�5�/e:��ܶ㗷¢�R�f�kzr;,�ti�<s({h���6��z�����¢m;��4R���f�׸���Ƒt��CQ1�$��\c2JE\���|ѩ�
�Tyb��G�� ~h_W�Gu�

�U~����i/��s����>Q��{Λ��}�1j�X�[��	Tj��W�f� �>�$=S>l��Kd�]\g)#�\��&6Aq�!���B��>�j$�2��g��VZz��-_n�j�A���N��m¾̏��"��,\+�'N��,t\<��"Z�h��Q�b5�Ѥ�=E�/��	�W���7b�a�9j�n�PM�۹�����5���MK�C��1,Fx
��'��"�^�.��|�{
�$LoE�G� |��~�+�>�"��_�N^�e]�D����-�D!�ͣ�f��(i���oA)l������k��)X�^}�FЈ�bHsc Y7���r�y��׍����D��J,U@����k�A��=�7'�c�8jNv~T�,������MsU1�A$��Ǣ�{-q�N���iʘ��|�D��6�h��ÝɫX�/p<���Ģq#6Rj��A(B|�"Dz$�`\x�e��7�I�A��l_����l�'uD���=�
�Y#(&�v>��jb����	�[$ !.��r��G�ʍ��� S�G��Lr���V� ��X��A�ӏ>4L�e����v��A��y.�_r�~3U����JR�y��e
 HL�@�3�U��S-lp�,H6�Il��QB=|�ICË�"��Ul�����<J�gl��A�4����m#�KL�D���G������/XsI=`����������YdFK@�wYȎ'&�O�I$���=��P� �K�E3����9����p��u�\t�)@��?ͧ���z�c��)��<�3S��B��k )�?��R�2���}.;iX=�9�[�7xK��E{S؀��c�Y��yK��]��M�$E�<Y���öi4:Bf`���	%ao�E���:�/-����3?p����䉈�>MH�1::H����S�\��d����V�)��.��ϖz�1�8?�U�J������U������,�mSd���e�'�]A7��'K�߃��lH^��cTHY!z��R���!�o�����]~gM�=��n,��ڙ&Py�5��i�}ZyQ$��=���򜯟4�og�Pa����^F�72_V?}�{����"gY>.\��M��W_F��	s���}ny�v�}�7�J���|���%\���n��f*D8����^�ռ��**������?l�Fꌫ ��q�������R�h��ZilŦJȌ�|� �Ҡ�s�����U@��77�98�T\��c��C�CY����ޑ�&������`�㠂�#F�l�~�'O['�����k����,NQC��_�p!����IiK#\-�C!l �a,�B)T`�j�l�7��i䡓�K��nطq�%r�h#+��)1��w-����6�Y,��-�Q{��~�|͔��`3�;F
^��Y��}�+�}lg�N�T���D}}=W�^9��J|�H��"7�Rj"Σ~�u���͢+*;E��m�#ˍ�+)�:I#TX��Hm��`������%��l�k�11�4��y){sf�﫚��$پP���
�`�`V��(-~��#J0�yf����M*4b� X\K���y3�QE�s�b��]Ź�V��^"����Gj���sj�v�iRR�Bp;��t4u����yX?"�	�Z���&ͮ�MN�r>����a��7�8�������Qb��E�A�"l��̔�
���6��퇔f�����.�e��D�h��?�������ؑ�����jG~��r2]���^��7JBzۍvs�z�,B��K{�:�
�`0Q���x��[S�Z�1����/�pu鵄���2�,ڍֹ4���KU��?����.�"+-:5����Z��V�����~`&����(�Tr�1�[�Y�!���7LOH������K�	� 	��2���G6g��R�)�e�|H��K�U�a�T
��&T!�pH�7�b���l#"|�q��3r"�3]��rr?�FŶ |����3�?.���`9���ȣ��o.'ΰAd�`w� �jl�l����w(�Z�)L�3R����s2�}���:��<��%H'3����gFW_�[~���i��i��e�x���
Q���}AKpT�T�� �-<\1
�Jܜ����iU��yZ�$B`a��jj�U0�����Xj�=0]��|���t��V���Rl�˘툷����̠N�}V�;mj��~�xϢo�8y��zQg������@RnZ��[`��߰��Cc�D�~�yDho�/�W,<W����S�؛����T���ƂM
"��pK/ys��>��P��˒�>��yCtK���x�u�p,d�&%�R�ՅBh�4w.�^/L�)h�v�u�N�|498�Ne�fiS	P�L�K'qE�"�;������_���7_Gv��iE(�8/�4����lX���Սͭ�l�
��=(V����ޓǃ��`q�;�w��yqZJ����ˎ�ز�[�>�ݦ�R�Ul�T�h8�Ti\c����.+�)l���(E�)X��"�,�X��KQ1�8d��'�,5�eꚸb[ce��x�$�B3?����"��d�+F"�c^ę"��S\,�0���}�AF�+f��j�i���la,2��-�'.T5L�]Deh9R޷��M�����0yu��9���x�D�A+��+�Y1P�|��pA�W�@.c��8�q˄\��PV�l?>%\�B4���u�σl�?�.e���Z���`{��'����VI�?����+_N�V�Z��R4a,q����ZN�o >"E�tU~I����%����^V
BU��+r!K�ZfG刌�dX�I ��e��6�0�{�����P/�G:uu�K8��c��-U5��p�b��Ɠ�_�؟�/��g�p��|M# ��.2PB�`�ĢB0X�DT�'�
y�j]��$�4n��f�p��ɟ�Sv�)��4Z;��5O^)�ɽ34�{�Na0���-��e�2c%Ag��z g�1���m�n)vt�����$?��$!�͍�_n����{�|�k'sy�� �WטyB�5��4�Å�����=�����_B�=��T��ބ�\�
�q���}wBn<(���~C������Г4����86I`�R��+~�)��ur�-�lb�B��c��)KW�R&C���KU��6��M@�Qѳ�V$m�`�X��\ ��4*K�>�P�����I������С
/�k�$�cR!�`�y23H�.�1��H3},�1�d�J�Y��������P_�I1ZFg+���^�L� Tպe�.��'c�c1��gT�BL��Ի$K��'� q��Zh	װ�,�f�B�L��t�h9E �#�(��C�m�l˛	%ɚ�K��M���B~�T�X�iXT1�V%V�E���M��-F��Gw;3�v��ռ���L�T�z_!1�"�]{
>�|y����1����()N,Cq>P^5�*ಹ�~����,|�%+E�L��0��/S�k�x�����j!!���9{׏6�7���$;�7%i���뾎�.������M��O�ĺ�3:�}�� ���o�~,���g�&����g~z#$����h�:�f"�p�"Q�w4n�9�GVД�U�� �B#Y���Ц��B���DH�����y�j���<ޟ�*O��C�gд�(�e�����4-䄀��%Y��b��ٵ�>�+���U�!Sq#a��$@eyMF�؄��~]�}]�s)rY����qz  ���y`�BS���ıHM3^Sk�kv� �-�pi'�5��C:/T�3q�}k�i�Dg�})C�ﵪ�� f<U��|ܨ0��4sn���8K�R�JD�~2pc�°F�!Z�c���mO"���|�Zs,��tj����a���7sn}|�4�T.˽���
��$����j>��H!�.����e��"��\v-���!��;�L@˱R1�?���)۠D���$���ӳ=j1.!s��]��O�<���gi8\��B'�87�� �'��c�Ez�7X����gVV�Uf�/����1�%��jo|~�{-mۢH����J���?���^H��+��6�|�KƲP-�n��`�Т�7��&��k�3��I�J��Z�JsFy��b	Z�H���5����DP�(5�m��r��{��4Aq�0���_P^~��)�0�����=��D�K\�<�T;ɴ>YS$ �B���Ƃ��]���P�!0�I�QZ�@ (qVZ9E��%.Y�b�\�������\�8 �pݤ0]|iDIHk/A,Z�q�K��8r� I�+�&���3*�qRSZ�ߡ�����w@Kī���N���+S���N.��ٮ� >~�5@��������oVΧ�M�[�ʲ�3��ߨkن�-�����yDН�N��`�p�MR�c��L[=S�)��wg��y�П�@�ܧihT2�b3������������#�U﨤��>���R�f�H�Z�e!g���%�NI����,��m��'��4��>���I�~|��]زD뭱�I�<dsE�骦�Ԥ����vb��r��Q���J���y���*�"\�w��>b@�*_>��6� f�¹�6po�q�G��:J��]t8���P�Ӎ�8�;HjǙ�RS2&���""&��Ch�B]�TgNd����(���%궑||�m��U)� �����v�7o ЅSD��+e"/�q�s�*	�C|�w���ɫ�ĳ'�e� 0�<����ާ��?�^t6Y����(X(�F��☔YL��n*�A?\�������SqOMlv���Ր��SL,ح>Y0mV5���~�EA����@�$@�,+���!�^<%�+</?���N�o��S�⊫_�Yq�{Z�[��jǃ�j*����ǨtS*_����pŌ��9��G�:�>d��w�Lȯ�:� ��7�W�D@����M�r�����>�/*���EIί��$�
��3����{�M�;ן�� ���,��f׀u��UT���� K~�� �iJ� 0=�!��%0�C��!@��ȃ[;XU�wU�7k�J�u��-�	\�x�=nS8L�>�^�_]>	���F�^��Q����E��2-1ۊFW��"�	'Gq�G��l�RXW<x��$�{�R���n���
&��޵Z����Y�[������A�gPk�So����c�Uhm1S��8,LK��b���TG�A�V��R�����$S#��s���<��u]W��	���2Ao���i��7��̋(�2jZY=����m��M��DW����������:�K��	���SPdc��]]�Q@E� c��7�l<bm�d�<�l��3HG��p�����aF,��)�2%>D�̆�c�)�'�Ip��:/�G�Mk%G�C'��K <Z%inpR���J��� D�;d O����Ah9Ds5 _�B#�꒽��o/@�!���~�Y~h�f$ڶ�:���}H8�i_��0�ID�ZC����pE�t\�8���b�e�q}Ē¹NZW���ER��df�[��+Cr�4��7zBf3�	|{�0����:j�t�P6���j߲�7J�$���Y�Mr=t��*n��B;�g���ڊ�N���䘺I�)?�vՠ���Q�M���	�5�-��YӜA�{��y�躦�����'�	�)������q��B߻H�(���z����k�k���*aW����`�����uZ�*���k����+j�xپ�@��v�����u��^|Ö��@Q��x�h�����E�/(%��#�fg��'ǘ�Y�g~��� >U6^{���R:ϱ����lkt�+-�n�z
2��#�� �j���A+>Z��tN"Ǝ�xt&��|��Ϣ��8H��1�b�p'w5j[g\�3p����:������]�ɣ�ʨ��qQ2J=�����(��[)w���1'��٪bX%&�m�7H�ʀ�=���)&���s���D�^�f,{�f��;҇!C-���\7��k"q ��gC4��� �"Io���v���D���bݸ�*���'���xB1��@e�Uo���|i627y4�C�E��\� ,�5�F� �6�Ja�,�VN9��S$)=� �G8�,��js��^}N-�P�B����E�h�}!�^�hKd��V�f��=N����"E�4��?�=��tG�2Q��a�2H�lBq���q��.~����6w����{7Y����[�P�r[�}�{�1�����	9��Ǥ���g�+�Fp���p��F�t�м�$�sڗ�{����t�'{�u]�����"�7?��`�H�f�l�ɼן6������8+����3�Dg�W0o�xPV{��ѣ=�8~%�*O�T)���N�����B��>�K~���&��{c�s�?�/&hJM�N	��?��"��&��f�O�Hs�G��V
��0�'����;��'��`�Ց~�`��M�[�[~~V�+��#g f�1%O/:Hg�o�e���y.n 8��e���ͻ���ǳ8�����cZ���Rj	b�X~���&�A�>yv ��&Idg��G�1��;�"�PVO���j�P��A�x.1�fZ�m�Q��� :&9�V%@��\���c1��d>�FQ��|k�p��XM�\����*��9���Z���n�#�}��"=_s8D��\�^�t8(&���4��o�<Z|f�w��Z$i�YCyҋ�~m�{�s�3H�ŭ�Dխ��#�����ۉoD�E��:Zy.��d�8ɋ�p��D
0hxP��?r��v��L��?�|�PCR�������@f��G�V8 ��RLr-�&��m.[m�`�d��W^��%�X����#�v��������Nfe�sR��9P����-N�z3�X���\"V�9&��C��k��b���xP\lJr�dߖΊB��2��S����zCN�r�yr�E�f����m�Y��-�_Bc�9�xw���=�k~ـ6 6,U�0�ʶG�_ؿg��
��3)K@C˽%v��Ee�G�h������C��l�o$p�z�p{�<�Ũ�?"����pSP�N�s���F��iۙ�ٵ��=n �yKځ���5�9��n-�)��쏁�t�1��j[ζ�\_�dC��Ǽ:��>s\C@���7��Og�2L�?�8�T������jr��ĝ�mr0��~��
\n"�r8l�$m$�g�婈�:ɜ�8SRDC*�;Y� ����r�H��C�%����%1�s.�� U�S�We�$ƽYkqb�A��q���LB }��瑈&#�R`l2/astn�ɷ#��7��Ld�B����jY-�5�������V��̷��jrܟLh5'�'E@r.4v I1T�n���B|�� d�C{m��Z�x}��M I����\2�T�n�S��"�\���4y*�4l/M�n��`���q��}bo��l�d�&$s
��t��$s=�?n�]�PZd݅-�W$\��r�#��r�Ҋg�yS��V�1j�t�ju1��W���}�C!��P��?�����/�r�E���������h�S@��]F��c����j ���A�rF�X^3)s`j�0�I9��Ɂ�����/�}���f�ģ$`�I��Z�u��t��s�hBc��!������|�6T3����J�Lj���
���#}�V�E*Unƨp���-x��L{F�bb,�zQ'�CN\u�)���I��^u��.Ey�Kk��ϠyZ��!
�,����U�ep`Q�o�G�1�f���v%r�A�:��	Z��E ���,LƻIE���j^�L���k1���`9�+��C�w�'�1d�bU�����w�leek|&ѹ���i=�Q�aU>��S+��W�3@#�GS�~s^5�"�
�L6��S8|Z.�j�7�X���w���5[X�Ej�[�;����������>�y��c(��w��� #��֙�UG��-����4�[�&. ��p��QIߠ5�L�6����dZ>_R�N����B:����g4X~cx�U�@����]�ejz��R%l�#�^o�_D��U����E���=MQt9�eY	�eN>m��-�h�IK�-��ۦRm��*m�I��/�ȸnc�آ �i�!�p�Jq{�|t�/W�M�����Z��/F�y�����QWd�|���'FѦJ����)q1Ri��G��O\	eIJJ��|��!2D���'/Q�T:8B��$J�cF������Oˮ��t�Ϯ`�v�_lǻy�V{{�#2ר���+�n,sl[.���^'���e��B�&��[J�`�P!3?�-9����3����b�C����ڟ�D��<N$�9�o
}�� �Ǫ�j"�����,h�R�	��̊d�T�I�'2y"���A'd��k�p��e6�Q�][��L=Đ#A(�:��!�׾��~|�r�h���doė�{���
ķ̣P�_*h(������ޅ���C�O2{q�H>@d���ŋ���(�<Y���ҏ���V����7� .���U��%ZI=�vy�����j�B�#��^�_t�Z_�e)��o��_�:�\qJٷ�?^qH�������ИbYn;}Y��>�I�����;����זV7�,����V)jp
���QA��@���5�Y �qM��� Iڨ�s� �T5"-�.Y]�d4��/4�B��˓x|��4�����u��d�7UC�µZC��H_� 
H�n���K6W%c5U�|��/X$�=�?��B�Hh��������&%�I���U��K����5��9])n.gR��L�[����zdEcÿ��5���@T���ag���ͳ���w0hx��C`�46�����b��E�2T	���>X'�X��BKIH-9#֞�x.�U�v|�'�~Br�oZ������	�И� (���M'�^�	Dc{�Ɇ�����TeD�rI��	B��g��e���q�Z��]��}I�h��#�wF!�2�JZ4��jg���1��N����Od�w���a���I2Ԑ�������x]�z4�(��{hv���7����ei�2���s?�Ȑ��(~�����F�>�0u�چ�K�I#Ix���S^��j}�L���mSw�#�?$J�pA�P(���k�:�8�p�9���Ѧ�"�$�;�;N�J�r��R�ǯ�t�:�����Oj}��(��8rK���:�b���:��V`{a��0��z��� j<�0z����g�|T4^ 爣���ă���^��_jVl�A5��_LDQ�S)��xt����b� �¸��)a!��](u���r�($_�9��#�j;=T"���<<�-��}0�V�w��Q����uC��M��2�~
���R�?�=�`�5��K:Dl�m��l���3$�����]��uT����+�U��"(k�������|�����-�:S�H[}�e��T�wd��8�r�+;8P?C	��E�Za�$U��P-�@�i�S���[7\��ʃ��]���P�9nQ0�"���b�l؁��Ď3�Hɱ�����f i�B_�C��/Z�-V��c�6ԝy򇿕�!���,�Q�
Ul!�r3v�6k�������<��?�J\<��"��Æ���Kُqq 6��C
R��q>ܜvaA�=�?(_��z��R�Ǿ�=
�Z��G��c;�#�t�u1��'�:�[当B�/vr�9�ӻ}
�EǶ�@zkI��1�?TEE눬�i"n�6g��=[���?��7||m",�c�`�Oul!^�q�ӕ�RU�g��Bȼ��X��7AD�dޮV���h@��;�9������jvZ-V����t'��e�Р�H{G���ǿ3y"@Z�;�+�|~�v@N��p�+�G�;�~�}F��E�HO�*�����J�I�Q������}5�\����v���D�s <�����FXv��1�2��:%T��V��?�I1��4�_�.�u׫�-�$�M	U᪀ŢGF^m_��e�N�V��ƭ8'��!
��?hA��v��޸Eݿ���4G� �KK��►ﵾw9����dL�V��#A��-)Z��T��տ��S	2s��C�Aj�@�NAm�h7���q#!�C6��Ia����8���z�-��nB���v_��'��)'3�_B[����G+I�����*[���A��)H5)������k�YYS��|�>�ϟ��8Xk��!�]]�t#�塔�-A�j���A�%��8ڃ��ҟ�5[do޼X��g�7'�ٱM���R@��@�`�]�@��`���Px����� ���Q_�k�#�\����C�=w9nه�W��D���>ݝ��4��ٕ����C⿟;@�a�(v��^ IC��NB:�=���������Gm����8s��yG�@�5B�T��4{aS�Q�����KNo�	��2�L=�Et[-�c1���l珙� �((�+`����*�-B䂜c>5aN*M>�Ar�B�~W��*7�z1����3=��9�a}��t/���f�U3�m�X�����D$���!iYqK�+��l�܏��zZ!2��ͻ���K��%�)f7�A������FJ�5|�������!7��w&�U�U��'�Bѯra��`_�y�c��z��@H
��v��S�ωƈ�h�!�1f��3�T)�R��$�_B
�3�[�1ԑ;�"hK���?(��=�x�UCE�ޞ�ە�c�����dB�S)Zb�=�/���n��K�m$ԭ�s�ą\��׽ `���"���XC�3�~�Nt�W�A�������B]��	�
7�b����[lƆ;�A�6\Ê���/~E���t��E<���!d���������'l߻]��H�Y�^���+h!>�F�J�/���^��q'�y�T�	�e�2
r���FAK���CSoi�$h�M���!�������-A����ٲq�:d���2�vV]{��_��W���ԉ+�{B/q7*��~飘��O3;��="�2O�{	����I�_o�-W�ˈ�z
�B��⊑�w$�!H5Ew��(�^�{�A�]X�QqG�����06�"�܅���b���a��@ݼފ 3��`������a�|��*&8�C�~�����j{��_/�"@���/�#��m)RνI�V�uC�f�yN}W��k�k������c-��	h��]S�`�Ę�]Va(����)]�u�q��&�������=?����̝GBJ�q���Yâ���
�f�X���0�QEVm��$����Q�/����Ճ>����������W��[�}������MbʂX��{n慽�C�ZNd45�_�:ن�	�6hW�k��b�	���g�Z�Q�l,���Lj\��'I��}�ܗ�:fn0�'U���jE�#q_�5e~F$xUM#% �C�h.85k�O@��q��L��Iݏ�����Mu&xD���==H�:���
| �
�\nTx�ЭS�f
A����!g�������#��a�X8!>�b�u���)f{�{>o҄ЅF�o�Uɛ�iH�9�lk[������n�oY�7z������9N4�UQ�]]�._�����{�%�3󏂱�J�Km��3�g�$|�mK���u!�񜟞�Ք�>2Qk}�Q��m�K˞�o��L��s=�r�8��7�c � ��(�!ؿ �XH!@\��9D.�����[�E�u��3C3��CJ����� -�� ���" CH#���twH7H�4H�t���y����}~��sű�c�}�}��2h���*(�:�����iI��]��������_P�0^���iѕR�L�T iL��c�0��L,���_Ū�z�ԕ���|��H@�L�QU�V�j����x��:2+@������Y/x��=�����N Ï��Ǐ$ׄr��y��+�9���Z�������j�D�KI*
ɔ%����]�?�R�K+�?�8�+�z@�ws7^}���*�J���� ��Đ�A1>���x����R�[ga@K|��xB�vI�P��z�Z�w�E���^�����s@JE�y�A�l{�y���L�`�q���d5���(��C��`�__�i�}Y��*U�6��7F�H9��[y{���������4�[���ʑX�[F/zw�g�i=Z��f�.�OܭD�*V�-:�y�~��oa��-�Vg���[U�" ?%�׫��wg�~�a�n�ݎz��EH�P&�p��z��Qr�S��r��|W2���U��-���Z��HFC�#��x��k1r�F�z�
��PAA>g'�ݰ]]���U������ё&�縆l$o4-�BV����s5~��	�����WWP�w���A�]lĪ�h6��w��n���yS5y���ª�	��Z�������zQA�x^���n�w��r�_ !.R3��h{"!>��M��RI� N���~�z��'˦����EY����ъ[m�P���r\[zT.ʗފ��R�w;"um�2�D�Ô|*豅S��]��y<ʖK`q�֕���	+C�d�뗒(Puq�������ߓޙ��P�89J�#�"��u��l���.1
~ȥm�{�ۦ����]�Sݚ�	����PQ ֈ�CH �U~
�yy�V������ݿ����ʌ��̚#r;d���>n�BB�(_/{���l��:�o�y��}nZ�>u3�!����"�������D����Mj�j��[Y����N,W���.�t2��/=��e�6��}B߼���V!���J��h;���sc��~��D�ࢊ�*��K���7��˨-�F����A�&,,:;��5~�������w� ��|dn�ݞz���:��yl MZ�3�G�A�ٸ�34s�L����pZ��*q��|�J��vn�x��f2��L��]-�(W�6E�"ۿ�v6���&b�c�C�� $&���^DE�8Y��
B�찋��Iׁ�f���� *�{e��g�:��V����%�MO��X��g���"�l�M�	��A�����ү�J�YT�=@��������0���xB�"L�G�^n��`n�w��{Է�
?2��UT`+G�X A*�R����� �����2���A<���z3`21�a���+U��&L�e�e0��X߱`p@����$I�Y��9ڕ�N��L �.;>�C��pӰ��2c����Fk��K4N�o��3$����S�&�,:�\���K^WU�5�AL�z�8�|$�<oN��]E�=�ޑ!�~�!��p���,��H�T6���	��yE�bD�ʉ�;�2�ۮR�����\��5gQ9��&��1����� ��2P��`��d��9�����ͣS�ôI��Q�D���
��/�e�='���;%4��2֘`���S=.�pR�	A\�{����;����x�4q��843�V�4�G� ���*I�gr�) �Y'l���`��_� <��"�w�`�{�%"��-����?g��B�os��Zu)-�q^t�P�9�$�|3�Is� �V����Ͽ�y���Qת�����e�VF��S��PO��fk��#��d"��;��Ä��+)�� &��e�}�9^0,�}�{fm��4�>�ג*�qV��rA^�+�R�{��~�uK����.�a�q����W��a��3D�> �?�pBr!��u'﷣}���!��n�GOL�uW�V:r�
��Ez�N�J�NkF��̸,ќe�+��P0��!p��;�d�.���,���(wN���W���]�	CD�[�܄�L�_xh��&�W|�k�7���ϑ��.>�΅�~���%p�L\<��7�Z��
�2�YaZڙ���B�&���'a};�WL�3���]?� �s_��������Y�q�Y��$��8��B.d�FO-��9�H�v�y��Z+�#K>�}�{)d	����Λbͪ*�f����g���m�Q)
��av%�I�=�{���r�yE�W���g�wț6`(N���/�����_��H|VL+Z �Gf����/�|�Rr�@;6]X����-���з�h�G���h���l�
�X��\�&��O���8��.���+��P a�o��'z�N���rr�»�b3n���7>~\S����1�tVs�jp�N�����@�vb���BAq�D�IbZYP�<м�#�]L�)GF�>P߁=x"�_6��EQ�te$`&��2�ُ;K/�m��l��j�̀���v�wf_6m�?�n�G�|�<�eVЎBEDꝗ�>��e[T��*����('���4�UT"OIIv#�X����˟ �PCgrwCr����H}pj6��Ʃ�l����>Iz���9r���X*�����%}�2yDu��d�܋�N���=��W
;��I��SU00X���S���cG���&��0x3(���Hǲ��j��u(����R�IO�U�s�t;a��WS�K�_(�y��Z�f"�[6�-���G���Zuh�]ϖ�t��vY���@R�J�l�s$`P��,;,n���{�do�h"�4"Q��GY.>K*�i�|Aطc0�%�b����E 2��MdS�K�&R����$�\BMD�K�H��0�e�FX������U%�@��T�Ah;:�7ao�N ̤�&� ��$Ip�h}��`�Wj�> f�&G���O���,9)��l;z����$W�m����k�T0ڞ@��;�I���z%}�����C�»�7�J3~�&vAY��I����F�؎�F��D���	����Cp���!����:�Ϛ��m��5��Vg��%jaT~��x���H�r5�}�zc�����jyb����i�v�+~U�$�M���ö�u����������[++��.`�k�����"�@�y?$X	{�Z��#e�hN��U�J���~v��Y����y�0���i�G�N��8��v���9�i�h�Q�`0a��GLc�^����4�a�G�#p�@XIW���:p�1�jSl:�}�8ο�9W���3^<��Gd����(�CM����#�k8���5�F�����+©���s+3�}� ��Cq-Wu��X�1QԼW����O� x60�������q���/�jx�Q{��F���K񄟨��+�.�Y����V�B����H��_�䛋p3t��Р���1�?�o⣏�.�W���M~/��~U���j}��L.5/\��v�˸�k6�[ێ�PW�:�����۷s�v"8�s:��m���濰�iP�"7%��N�~n�|�a'"������žh��l$Ā}[��� ��/� @H����Bۡ�gG�!k��Ԧ+�x����Sq���^�ӓ����SHȫ>����M������V�hfg��Ue"�R_����)!*��X���`ߐ[�:��ۺ*[?�_��k���-���M��ݭ'���+�u&e;�Рͳ���#���Q��'AX�gV�<7:�ߑI��z����H[C�Y�����bV�[뻤1^A���r����*���H�����w���Ϫe� �1o��r���)�=�)�6b�f�e�H���k�}V�i�\۵
�dM��qC���ʷ���G5����i�hs����ǧ{����K�h�?��Bjk\��O��Z�d�z���h,��6h./�[��EG=���r��_���oNl!�cۊ2��a���W��x�L���L;�[�+~�z��NU�)v'y��.F�៕��@7S7���RG�4	��3\JlƧ��ރ��W�C�h��t���&<"�Ѥ=���΢C0�P!<��jk�#�����rDZ�#Hf E�[� T���������� �>��x6�Q�e��i��w���A.�z@�霾õVʖL?����l�tN��+����4&�Qo��5Fj�'���1�BInJ2�')�^��i���v�1
T,+�u��R�$s�=�ɻ��#�0W�KB_aQJB4��������ӬO���(����6b���� ���ĉ��7�G�Hࣿ:�⣢�/M�⃒T�tTB�����֖�Ԝ /
���/�2���J��L�נۺ(Z(WW�|�D�����W�?�Ǘ�cM��dC��6x]��A���9k#/�P���]�A�*�U�/GI��b=�g�a<u��UBBq��f�S�؃�5ġ*�^ �!�Bu�"���>u�\WU�ž̧^L-A�M"�"�O�}&��`㇙��[ъ�v���Ҷs�g�0�'fA?��Q
a�ĳ��������*z�sz�.�{�����aR>�x�����H}j���8XY ��Sg\kc|���h5����>�����eq3f���l��N��k�'�tE��wI�Z �\�#A6��T_ˀ� l�%Ƅ�#�h̓� ����DS"����T���@�'P�F�"�i{����=�����"%����O��1��y7u�ܭ^Î*3~g�÷�ѯ�4>��B��'b�r/3�0�!���bXڳâ�Uy@�7߻����	x�i�2zm%C�� O�,���r�;7�9�܆�r�:_k�o�Xк�6[�3ة�Y��F<���A��k�w�(��C����|�������.CK�<���w!��u�*6a�c������{�����7��q���<=�5��>z�9�)��s7F��a�Ϡu�)N�"T�ݍ�.&"�8a��XC�{����e����++��"�rN�7��K}������"��<?&��%��}۾�>���mG̀B]�{-��׮�T�11n-O��P���wX��_q��߃A�Xk��f�[�=y��j��gR�aROv����wU>ܟ���yg��&CO=�z�������Rf�4����.�0�R^٬�~�A�DqM9�k7r@4<cQ�8�e�v�;�_`CL���"IA�%��2Y>�	h2�`�V�ґ_�P��xOI#�5��Qߗl
}r>���隣ǮM#�p-�SA���?ao�5�㫉�s^\dܡ�	���?Έ0_������02���?��ݏ}����e2�Gu�spV��ٔ�	�Y������.߾�Qz�z�sY�(��( ]�=)B����W�K۠��6�oz����X/�:�8�x�KK7o�c���)�˝_k������_Ad��=3g�L-�VϪ�5w]�L�C���x�|hu0w�1i�h�R��e��R�4���N�8�-�g�*�fKe�g=��[ �*���ۙ��'��������f������8j�Ϸı*=�A�҈C"�g�<)�#�#M�Œ�3���GE+�/���XCMV](�iD���Q^��w���yK��ѳ�{�>o��g{�%M��'X��N�E��c�$��/�%tn�A+�/������q�߮��:Tq󕂰"r$M�o�4�еRu��Շ����8xˍ]dH��w0��S돵��%xBU|���w'����٠��+}�TKT=:�~j�k�Z�3��g�#8Jq��:��	��5�5 ��K[���Gm۱­A}_ɩ;�F����Ӈ��e �����?��0W�~K":0�T��Mؾ�ה����;� ;�L��"�ɫb��RbS�m��e�D�'ݫm��ѱ��L%��O靋^�%���#qO�~���^���x�R�
ۢ��L���<|R�A'ۙ���7��9\���6�����0`��G)����d�*������6��Em���\��e�E���f���rU�9'��m{ڻy���=�6Y]��D����h\� �F*XNl��r�����h�؈����u���8�e5~f���4;��Ξ&�gNEj&�tƱvols������̶��veJ^n����N?�rss���[D+�rb��p�tU���,7ե����y�'��-���Y�F�k3I�+g�4e+#:�bܳ,=��C�{-=�&ʁC�c�aG�h�U���F�i*՝��k
�B[��� J�ta�5�A�=%.����Jv�#�Y�x�����u�W�])����Jŝˊ�M�(??�d�[�c)���8ܶ�]��/~�^hFͅ����n��Jկ����)�T��Ʋ����zf������*��@��?H��Y�d&=��+UK��eA@p� �"�sZ��q䓌ݠ^V�[)6A�"��3ѻe���c�O�dt<���,Kg��f6CuM��#���o��N�>�[����;�-\�ƒ�d5C�����c�ق؇���G�vδ���������tW�\w����
"��Z�Xd�s��)E}�=��H1U֫�}�r"���z�C����UƸ�>Z'r�@͇J7l���v��Y@�CL������\��~���k�ŀ.�ρF�A�����Ĳ�ں9�PWi�� Cȇ��L�^�d:=i����"�������B�۔O\.����DV�_��!�r��Y�ŝ
�{̗P{C��n�~B�o�>pq���h�L;z ǒŇô1�)���A��Й�>S�6Y�_n�e���ad��j������w�	�>����3-D{���;Р��̸Pכd�Yg��K5����Ĳn�(��״�����:��H�1�5�SP������W����r���`�Du��6��T���v�}mnm=�������:����3`�J��BJh)n� T�{����j�3�4�w�I�?�&�v�+�7��m�MO���4#S��6�wfk��H���Xʭ��?�Q`%�Ki 6��*����3����t�����SvݢE��F�U��^M�-�x�\q��)#�� ���9Q!k-�T�^�.�r"w�}�}�5uw��ͦ�]+ gdR�{��ij=O��7��!�f�0�?�v����U��O��h�:�p�־�mS�Wh�@!�j�G��u+N���G	�)��|���s�$����-}��G��V�2}��x�|ŕ�� }�0GPe�C܉�?���F�TS"���
��<�#�i����P�B��J�<�M}V�F�sBՀ3�8��4�٢�ï���|��ʠ2����s/=l�d!�_���������(�>c��
_�A��WT���jL`b2l���2�����Ҏ��@茙F¬,sݦ.�m�^��/%-�H��;n�j���Aw6�Q���/�κJm���6~�oZ�z6�aY��\
{�r�ZH��N��m��І��0����3�׵7aѳS�^�'�#�K�O���6�8�� Z�"����
����T����`Gf�dĽ�¨tː�g
�{m�zO5��w��m>�Oy���߻)MĩsjӋ������*B����߼}+e�}��@E�Є��[�OA�wq�����X��1�
�|�T��v5pj\��m0i���ǂ�]� �%�����5�?��o����>���B�l.����o*#�iq<���ذ�y��W��E"��i����".�]f~��?X������z�b9��*}�a�J���R,���y��}��e��q��]hÔ�<	>:N��=�QP��".�|�J��.�\Yf���Y� ��ϳ���3%T������
8�.j9��f���3�-��@�<���3 ����>at����9=E��l�[5Y>�����w���+s��N�n0��E�3�X0�͵�v�"�0A�<����zQ�)N[q���н���ޥ�G�����A���
���S�x;�A���%>#ipW�8H(à(-�޹;#!}���ȷe]����=��T��Wo��m�k;���G+m2��w�y��>3�s�N�Zc*5_��QUK�*�x,��#lG�`�ފ^ԉ��!�$���@&\��K��9��'I�զ*;R��4)�dS�G{g��7&�o��9#h����Z1�J����H�ɭ��-U��7�!��,?ws�n�����K��2���lq�(i̯3��I��e�w��y�ա�F=�Q�hv]pV���t�}����Ĭ���w�O�ū;[ɱIP&ڶ�l�P-巸,羞$@�C�;2����%pu�|:��.�rs	b Z�g C�M�qvH���0텱(Օ@+ 1r�*�<wl��Z�nZ4o9�~W�t�{Z�E�^�`�ǽ`�r���JWiLEb�G?�k����J}�8�w��{��w|:n�g{)��&1e�2�X}/$��ccI�3N3��%]�6����7����J�J�!����D���$�S\�����_p����34���u2��k�9Xj�))�#=��E�x9�?z�֣�㢛�#�}U��UG[��ӂ�q��WH����
|?��0%2���U����L�����;
33�
����ќ����=�ϳn����z  
a h~�h>�G6i�߲��X���:����h�{�������M��)v��6��Ք�����^O����%E�2gt[N��n��Ǽ��_c���TS4暂ã�%i=D{����{�����
d���n�O=��(�Ym���z��D7
��e��G����ȱ秅H�����z�iI���=pn������S��B�6�(��`p]f�P�G�.�$���!<��
Q��ٖ�>����vB{��O�C�����]!���Q��[җ��c��5M��~��3��7�{�:�,��]{���cJ>Qd�]�@���NXt�A��ᰇ��^���bg�u�3L�#m��a�T����M����Q�!٤oKv塿�n��)Z����7��d��QUY9�H\4�&�v{���+`�,����HĀot����q���5{4���a�u��Kϖ����k�㔋2�T����M;�-:����@j��MExG�j�E�[���T�-��Y� &�¡�oӘ�<7G�-d�'/<��؋��j�'#a]�r,��?z�a����9����8���J�.]AOn�2m��\�.��[�Kr�[r�ԛ@4�Xi����YV]�%���?�Fb���Zae��n%ݕ�CU���q�����Τt�B�v P����|n*����蕾�<�[?/��w����6nH��lC_�Q4�i_�����;���d�`����{"��j#������v��ࠝ8��8��\�n>�|�j^�|i;��p�P��r��hb��ajc�`�V��Yj��s�n�g��b���=��(Ä��}*{�����SGeͤ��9�9*���书h�y7��N�Sˣt�ej��q�oR3�{Y�5N�'��7�uXo��(��)��E9i�&W����.c˩v�?p����5��㕊�6�`!T�I�Aͺ��fs����'C4�����pzjj����x5)�Ͳ��;Gbj ��٨>�<@eDs��v��V�h��3�3$ΝΧ�S�
8�;��Z�JZ;;�y}���#}��Ɣ�n}'�Q��hu=zv���V���8wC�<�~5��"��7C��RA���p	Чr��m�I�aZF��]t�8
��?6�*U�����_�ބw_��K�y]��r�ΤXg���h����J�]wSY����1��s������s�8��*Ez������� .�-��ѤT�ʌ����tE�O��u^��%���=茑c�iJ���K����}��Q��Wg�ݾ����V�֝Aj3X��پ�;?Κ�$]	d��6�����O[�o�<1��lHr�%Tؔ�cW�,�����2::)	|��w����՟�*�b;�&�����X&���m�����6�uM��h �_s	��a����w܃���y���kr�9I�����8�+]�U�GH��wB��;c�E=��u0��n��Rd-'EN)�_t�r~~K2��r�X�m��Puýy���`��~�C-ڒ�	���ؚ�mH	�$�>�q_h��Sf}�k�|rc
9��q�(�ޢ�ݞӠ�K�>��TW{�@���Qo��D�W[Jl�C�<HE?1B1����,�܈�W=5��տ�T���N�M]����%`Äu����D�D|��O)�SS�+�+�����ߖE5�h�P�����3�M���I�ɻ��S��Qa�%��K��Cd�E��� �[�j2��>��Nr������X0榮���\����	�Λ���:�x��G%��u�ka&M_{t���.���@j��mLR�d�'?5�O>�0P���jd��替^v�c�7�6"������l��C����Q,y�Zf��*�*������wOoo��� Ἀ��>W�s	l����·���h���5�[�W����M.�
,\gû?L.�7�)�����	�����ݜK߹��=.Mq���
,�����N�2+t^w��;���p²"H�P�fL:ex�n��u�5��P�{~Coˮ�	RpR0����`,0������I��d�i�7X΁h3?
K���1�� ��t����6θc�y3NsҟI]w�O����8O��&OJ�6����"�Œ�HJ]���B)?��f8ƚ�%��ݦ��w�c�?�h}�r%���]�X�� [�0�ZN�p&�C��Ap��a?�b��R����Z��r�&�)�*U�[8��L$�K D�1kfh�J�0[�<h� �rT�?���� q�w����o�`6�N
��?�.[����q�_a�:�;��4EtMU��'u!Z�Ӹ���Rg�C4�j��^����bG�y�E�+���M�2|~�8���p^D�}�gJc�(w�1�vI'���2�<�O�_��]�3ƻ�*���4��6�}�S]��B�4�b�T�������6�g�
s#qy(0�N�����d<q?~�I�$���e�ѽ�	V�NqgC�m��{,��@�/�tRe)])�>�Bv�j%ITf�#I���D*���΂W����M�m�N0�X7�UM�9��Д0J�]G��@^�+V�t��^�tEE��*�.�{���j�#�1A�/�n�N['b�⡛��(C�B�)2G���ڿ~|!��9R�#�0����N(�<�Y4"��x�	�~䙼!
��mDλq	��ܞ�M��L�~n�����Xhm�8�#��rH�/��S]����uLj�{T���[�+O�v�b�@�q�����k�\�=o�@��>Z�� z������\���)��t��-��g
�� ,�]����w0�:fq`��>��7��y�Mn�}���T�{:��Ir�>��zE`y:L��RA��*�lZ���[I�Xb���t�3�5�Q����{d���T�y�����B'Z#6fsCS#şoɆM�D��
V����%6����pz�8����J��%�rR׾8\]N١�T��I�p>�؋���h�(7rD�zOm^�R/\NԤv���8���,�G	%��t�;����4Gj�;Ğ��ыйE�8�ǭN2��k��M&f�.��s���-�	�=��b� 0�\]OR>����1�!8��A��¡;e"����w���'��e�z�rG2�l�H�ݙ�u���\�|B"8��n����""����P
V 8�-$����l��vv���D���,�ٸ��ګtU�z	�
 Y�����d����a/���F~���3���7%>ե.,�/��"����|����ۆ�.��/a�̅�� �u%l�kM��~	mĞd�Dq�]LO[g:���VI���>̀~�
t.4>N�\5��<N�H�RuwMJ��y�E��6d�<,� �B���?߸R�e3r��0l__����}�i�/���}Ӆ�����^7�o�ˇ�K�ӷ�Q��+�-�8����	6���Cxb���tqW��j�w�����2�$�ǐ�ƂhfX�cn�{	��\1�f�uY�bH;,mĘ29�>̰�(�'*��W�}Vayp5����k���S�ll�5�xme|�$=NR���B���~%�^ga�
��%����#M����S�H�;<�ÂU�jiii�# )y���r�J{Fb}����,�U��o�5|�ht2s����Ts�	U�Fρa���4�&u�]{)&��1�p]��F�P�<�؍]#�]$��MaJ[m
?�\~��΋)�Z�)��<K\^�Vt�L��wƱH�HN&/�!����,@v#(��2�����!0�o���=@Q�\��,~Qӻ=zr7����nM���Zh;ݝ:Y}y����`ݰ)�q��%�r�R� �#����=��ȵ��U3��E�k��i���5����~r�%� �k�+ҫ�����r�٥�W2��ը�|�b�D����nA����l؋�NtF��b�w:��=�XO�l\y�����.f^�`�-�fܴ�n����89���X�����
�L���Z ��~��	��A(Q���A��~�)���,D�»��"��ϙ|I+�2`p����)�K��5��f��;���c��Å`��ǩ'���`�̺9M�Nl�����<%��C+j���A���A{w���$��+jg��  u$�e3lU�8�~)���^r�����v�	�<��D��F��D�d��������k0�O��A:����ӊG���%��jw�)��ttU����� (Y�`��ߣ�l(V(�j�����u���DzSx��R���.Rֺ	c$Ne�~Θ�fl�I�A4����LT8�%�p����)�������Rt�Ĥe䵳�«0�<WF�h��Av���PRd,�G��q����r)��I!�ۘ(x�pgn܃���3��'Z!�m������?��A82ɵ��/e����t�cfǜ�c���c��ͪP��XO�'i���ku>y�g��SX�Џ瞳�F�B@d�A�,W�ϝ��Z���zI��@$-�p/>w�8Gֶ.���?��u3��jB	x�±k�O�Á�n��P�{a�_H��!w��2��!��)t�2��*��|>ZM��4��~/[���ӰG���+�ۄ]�8v��4E�K=���, �����퍱ƛs�u���r#�>��
�<�1�5���`!�I�ٽ۔��
w|ff�	;�^�[S���y/������Şf?�L]�Gr�����HI-��p�Q�R(�Hr�ͮS��yÏ(n��ޮ�Q�\��l��Im�YR�%�k��F�S'��^�ӓxq���1���o�mcg�s�Iu7�
�[4������
�#�*�����~���&�il�����2����1� ���
)������[�a3%��@Q���@\�_f��6��:���io/?6��v|�PQ ��	 ���Kt�ϵ8�[��gC]�}ڥ��P[��zet��9p���TH�S�h�c�^�הy�㷐�L~�( �A���K������D'1*�;{Ǌq��{���1!,�;�箇��m��G�F�I��#�.�/]��מSK@m�������!ze0���q��$.*k�,+��VŃ.��7�<}�-�?��~@qaa-���J�@B0��_({�[�-����b��3�7B(�>aF��<(#��'��Ĝ+RO~^�W"ˠd�#�<��xEB%M���i��6Y��Vf����/e�<�4>ې���scz/{<�el�lƍP�|����O#��NÍ�aAe��Î5a�P�D�W���B>�w� ���Ng[nf�E@�31����:6��?�h���`�8IB|vՃ��d/�5N�
��X��TB���ӏ���D�6���H@dH�#	�?��l��O\>���trӍ�ʙ�N�����"b$=&��8(�H+j�[��7ڌdV��h ���<f^���yЈ���p��t����ȧ'++�t?=�[k%�ףN}�z[�ҷ\
�^'�����i������Qe��]�8I�I�Ȋ���������(߬*Bg�0��<z�]�*l(��!�Qp��ޗ^l��7���Q���\
�I5�7��1�;����o�T��~�k:����jRTH����()��R��AyC���M��k�1��,>(���|ӳ��!HM�O��J�fk��E��`�]d/.L*Ē��d����y���F��������J^�Ư+�,-��0k{�jd%����0��2��4�qYp!=���� 	��{G��#�QF�����s���_�X����$3?��Y�;p�X��QI�"#x�I,�&�6���)u6*$���>�^a��[��2"�!b5$��# �'��L�n;\vl��p� OC��-1c�B>�=oU,�c��� DER����[�r{)��~��n�ȐP\�m�b(BW�d������A�B��S�2I}3�\r�s���ѣ�K��3ަ'�)-u�6h��շ	���0+��S!��an��<���u�ρY��?_,�Wޟ1����v��>��缗}�/]�UǽY�����j8<�z|�����F��N�i�����ף�֛Z�+��ҿ5[ۍ��.�c!ΐ��m�"4=�s�(���ttZk�o�,�!1�u��/�@)7�U���@�����]2��#���2C���%H��̜�"[����4Y�{�[n�aU��5Y�2���^g+X'��I�p�Κ���a�*�} �k@%OQ/jd-2D�p�������j���Д�[($���7NPm�)��|�ʆ���SOtb���ү �Wv��+�����P�ḿN�w}r(��W���E(�]e�/��ζ" I�"����lg�N�ezC�~i�>zh"NaZ���p�<��KK�760�ɲi._����Çf1т�����eE�ߕl�)Y�BP�}��|٥���A�.��!,S��Ef; ʁ����[���7n����X���Co+=au������#����Ï�7W���x;�����t2���\�B��Я EgPf ���P���
HUkߙd�Ē�^|-���㕪7��D���� �~6�}��Yd�2��<AH��\ J��O�x�|k=Z��1�-ݶWg㼵B̖�M6,��v0�\���W�ov�i"2���O]����~�S��|���}բ)1hɕٵ���d��șx�w��,)B���	�Y_J�c�����=J�����wʼ��}� 5J�r�e��Gx��0ьQ��jM�X��E�b$5!���'�7���Y�����+�U|����`�eYQ�TǦ�1In24i�ӣ�2i�O�29��5\�0-S�e��rΈч:�T�x�*�76n�mV�.���(��KJ�@4��(CG��)ﺏY���{j/@vg^?Ss����hC�`���L�?y1�s���a�YJ@W�`��%�v&+͋9��&nx����1g�hg���Wp]R�{�6����ƅ����H�a���rO}�����1U)[�V�-�uK��3�ޡX4�]����� io$���G����׆(*s��4��@_��$i�q�/���X��A�-x�������O0�}DU�X3�d+*�h�{{�]|�<�z��s��A�D1`p0X;\I�(T��\�T��5����<%�!yS&7Q�po4�(�[r�0ٺ�zsY�)oH+��ĉ��Q��"fZ�@�+ԈC����3P��>vR^{58i�k�gyȶ�i�u�j#��@�(�tx�38n�����M����G{�sz�M��T.tOߨQep�<��b�%>�ߌ��@~�y:�P2����%��T�Xj�Ų��^��az��$c�|*��E�&�NO�+�r�b�,��[�H�ܫ�����8�᝔W�r�I.+�dC��׋;򧻷Ğ�Fb��;U&��Z'��3l�ܚ���%���N+�T��u6��w�_�O�G���X�n��zV	pͿ��,�4��8 �T.�S7^4=N��- �ⷣ.�;<%�CV��gt�&���Y%
�R����>�I�B���G����[�7���6F��GqF�I�L����A	�m��q>�Eb�����d]��$kD�l�;��@o�*&F^�
/�Q(��ɏd��bU�&ЧD�ʘ�i�+��a��$�q�C��0���n��.��1�}�1�o��mw_������β{I�-
P�$[Pq��XЕP E�b���g���
Ŗ
���}��ǈ�a�z���V$kѸ�d~
*�/��1"�VB)�-�S
��C��>�Qrk����EL���0�ɠ��=f�ųE�?���������N���I4���m�~�ғ")u�?� �~�f\�˫�܀�v�'��ӟ��G[��;_D���"�nw��?���:Hfίɽ,̶L�/>�z+m kǺ}1b�H5I��i�>8�{C�
izoU�'G u{Y�i���� ��U˧�a���"g���Q��Qm��3� (�!Hw�HI)��=tw8�(� ]#(C��RJ7�t�J�½�����2��9�y�~b�������ky�g�����1���s=��<)��q�/�HȽݬ��j�w�}ᇔ�Z�a��%<u,��6f��=x���e�0o�d�g9��$#--T��m��d��?kԷ�tw{��F)*��m��������J�[�*��$�x���<-�H�k���~���;q	`f32=噈��,E7J���P�C��o*�6��deT���w�2_�ל*�b��:��Y$���A��±K7-?���]� �_�{��i��8�U�'
?QA��Ȣ���<�Ξ����3��@L�U������É�v>R�e!yMm~sI����/ږ�-1�,du��%�����x��ȝ��tad3�8�C��D�g	O���BNg�z}��W��A�/U�}O- y�L�+���o���;��U������*���3`'IG�4j���̣c'�������Z)M��I��T�90����c����Y�Я����ŦIpǤ�-��B���	'B�� '��t�X�ϳ�o'��	�.6<F�4B�#��Ğ�ƒ�..A�n@����@U�/��M��(��H!�,���W����j�)@"�da��+������BaȈ���G�m��v�1[���:�����k�7%��������e
C+_�OLp�lO♣�B�w~i�A�WvB�F6�7Y�w�)^�R��N=B��˾i:w��dqB��̱��g]��OR!�gz�5�R}~:� 8(��[#p���ȶ��-:'P�PHդM����}��X��U��=���h9�FL'�៼j�����t��>���6G�T��C��`g����6�{�>>:��;��T��D\q<�&���t��p���2}�W�ET6��*,=Ӭ�ċ��B�=.�dЧ�B�������}�)ټD4�X/Oq����w��b�n�Z�G���7�p�;�g"K��;�9X�ꓬ�}M��N�e2��I�� _9טm��+x�L����h�*�(J)z�t(Y��y(Azʘ�a�i��;�P���0"/I�AЍ֍3'	Ǧ���^��N/��)@?[4��viɿ�hB��P}w�����iTn��'_?�f��l��$�GC�q��\����S��}�0`F��~:"��)m��h�Ѵ��P�:+���������[�� �.�FV&a?O��XҭKD�b~,�b�C��O� �+˯��L��Vn&����ۄL�S,�4><#�`���b�e����H5���]�w_\���$�X$���U�+�Sa�ʱ}�"��v'���ZMK����x�X|�,����tM���gG�=����蹈�1>��!�~Θˡ�E"��I|�j����`E�b�q U�c\g����l8�5�݉���U��gWj~�<��JPcǎ�}�Աt�����;�m�k�T�*����-z�*�Τ�7�s5�?�]|��B��J2�)��J<{�ɇ��67�X"n���p�(Y6k/$U�b�e�}��ApZ�%i�Ps�r��%s����l��<{2<�39 ,V�2?R�Xh��k�L�H�۟��d�������C>fh��Wr?��VG<%�|���2����X=xϸ�y�f��y�k���$^����LAW1K@�z��f�y��,�l���V5�[����N �k��LB>�Y��!s ����Z���.iJ��7��H�[�������ye�D���i-逈��Q ��u	G�����I����e���=����,^Id��?���{1hs5��S(?����@v{-���Pb�*q�~���LU{Ü���U(O��>\�L�b�q�C��A&�/T�fG/�AvW9��c���s�4�wi�0R+��ݒ�*�h���$bM����_Z�F�����$v𾸫а��0"7��ª1ӯ|"�P5Ԍ��?�t��Q�,�ޅk�!Г�b��z��Q+C���>Q�A�0@����x_�_ ��G �\b-c�o�E������!F����q��כx�4��π���@�\���{}�"#�O�y�w!�=&��b�:�\���~ �#}�4,�L7�Y�q����a�I%�i_��$�h�C��:#@Z�z�k�lM�m�m��>�����|��Z��Fh
·,=	���e>\0/�b��*c���-١5Q��:����(�[��u����Ur��_*�%zb_g��f+��Z�4�v��-����t@MmB�ԧ��S��uR�e�Ηh�(�(ݢf�]��=ɕ�/���D���:��~q�G�Z��3��0b��Hb �u��m��bQkAg^H�uJ�b�xҎL	湟9u�������g��C��W %^Uq<%�[�F �#�>�ȯ wI�����/v��o�e�|�7Ҹ���WU�� rd��0�:�1@RIj=��]]�C�xn��������j�}S�Z;�Vvg�dth��Ո'����h`�M(b��.���<Ƙ8�פּ^#��H���$��HԈ��9%P[���=��q�d�|�iv2���Au��w��A����O�:ߒ��>����P�� -ev�_Ƅ����\P�S�ٽci��ٯ�{�\h���Ӝ�����G:���1�G;h^����?fs���D��(�S� �+��--z@��й���� ʯd���]Y��r�#j�&��Veؒ2���W,�&����3�A�t}�����D�z��LFޟ�
f+%��i#lZ����^gq@i(�C�'����@��* ������4�On\C1�,-8^�G�#HCC,���7�K�e��3��g,�u5������7Օ�����-� ��;׊g�L�qRd٭��9�gC�/[����� ض��� u$B�! ܯ��T�@�%��8�E���&�&�@�JT٤��p�y���J^A{LV�8�ֱ1�4�� {���VEjf��]�u�Y` �$]�����݄Xy$����BV����ѭ��3�����)�r!�h�9���*�`%��<#�aK)ϴ��"Y����яj,��R|@����ΫWp�E�y_[P�Kj�}�7'�!��}�͕KJ�WDJ2*7V�5��[ߎN2��N1E����q��C}�����v"맲�H���Fm�k�ڃ��6Ɍ�+0B��n�F�Gb����ʠ���v��0L��e�G�
������o[>�O�rL�!2l��ѐ�9kMQ�mڻ�싏N.9`R���ٷӯ��'1��C�Eފr�e�l�~�o�N\��q���e]p�!W���p��ԚC�^?R'+��/��Dpxނj���DK)Ju?�F�:LT|�J抭.g׬�,�bd%/]g���R��;�*�ܗ|�Hk�	(��o��a~����9�q@�߰C��OKvm�`���M��^.%;dgڌ�z�̬m9Dy`!�t�;3���!B�O]��)5����� �hb��mz?�{�DV�zLi��!R0G ��5%$�@_$f�IΎ�^�T���wRuh��ɚ��l�ZKۧ�?K1\ܰ������jnu�umr�����I뚤a��a�Vh�,JṰ|�1}�1��5 ^|�σV���̚����^ܲ�}�[O����\*��X��H�z�_l��1lT��d�h%\"Tp�~9R��oL+t��gF�&������q��JpKȍ{=a�yj.�a�Ӏ�������� ��1�T^M�<���v��B6b��v� P�P+G� ϲX2�F:-�N�z�qr���9��	(�A*��o&�<&G���&N��f�f���1�-����o!�-ǐ��=���r��]\!���4]�Q-R�������v����h��K5;�������;��������!_w�3�e�0�'�s8��&�凪|L���c医D}�\_)L��s �u)Α����2<�0Dʗ?����Ն��?���g�S��ݓ����1 Q�YlP8T���sY|&&&��,!�L�hT(	B�������[c��ٿ�������m|�]|\����6�m[����.�� ����2ۯ��`��xNQnL��b����m��u& �_YQ��>�(��YӬG1{�6o_T:�Sml�:g��eF:f�k*X���������K�u+o#�S��y���v_�<�2{��\��"L�����OcϪ��Զ/��C�],S�ܲ]����w?��sX>�B`8�,�� 2�,7����ku�D���?���l#��A3�mGC۳��l���Y����FYo<��,˓�%X��ʰ��n��Y���<�T3"x`2!mf��\Q��o��U�-}w��H�nJa�ҡ�)�(N�m}�������SWH!0Q�\7{��%'.�ж�St(b�:��Nkf9��E��nm(+�kB������m�44��>idR�?�7.�
i87�k0���Ym3�����"��q��?ί��ȯw������:W���i���I�'#�>w4��D���j`a{U��P
{�2��K;O���Z/�Q�vgxp�tF��F��|ھ]g�~	�yc%��o9��'�l�^=W*�^��i�&x���i�;&.s	��������I:����jypF[[�9�jMvc��Gcf�?5�ˈۖE� ^Ik�_�$���F0��80���k�? _D����E݈���<���6�t��J���A2�T'������b�-���3�	���c�/S�^^������aX��@
Gl�?�`2y��娯���-qhRL�7=��{Ro)�h����%�/����p��+i�7��w�7��:��(���W�hZܙ�p�UUCwɼ�w��U_/7�5xQ�^��[��L�A�����L����}W>)����S���^�ea�=��%r~9x�*�*]��"�Ibx��E�����l��+��1�Q�j����ڸ��2t� �E�_�縀Z�1$_J65Mn�El�<��*�lι�)�0�9�~�֛�50�"X	׼�C����_<��"E�uwr̉f��-ђ�5��1�q�����C,�r�:��H��)�)�,���'t,�i*� ��M��2v}���}������qԿ�Q��E��ԣ�m��wq`��:��b�s�C����.��B�ON�d�Y���!�=M����g�5M�9������u<>��?F���;T�^@`̊P̖�$�h#�G�=��ꅮ�ɯ9~t�_6�����gy��6� "0N#��G����9���y60(�O�1)2�o0��[蘻y6d�o�UCrR�.d���Xj�����g�w�Y��z� �v�Ӈ%���������̂�AQ�z���u�P���X�����f7�|f��' ��[�$<�4%�\���]�:3��x� [��﷓�FoU��l�\��sp�����d��ɯ���N�Q�'��*܄�7���em��?��~G��v�9ޱU&��Y����
`�~u<u���%�W��ʎ�l?���߃�������q)ѐ����"A�R��̟;��r���#�3������Z���	,~E}*q]ٽ�G
.�����i�]�c���o|��R�gwY� ��x���H/&	ň�$͌y;:�Km�E�ڛ��~�� +(Y�e���i<t��+� ��, n"��$�j�ْߕ�@��Uud�f~��	C9~6����D%�6N!�%.fb6�D�y��Q`��u��>�����z1���wk��Y���:�������PFOBAƫյ4J���5�@�i�Q�D�C��hֲɜ�\(%g���Wiɍ�]i�g��;�r�.�Dj%�g#����ƔՒ$O��X�-��Gq+$9�#ƙ�8??��z�e)#�<��j�A���|��O��=ּ���'W^�j�8�z���=�E�������O~~�:�gf+�똘���#qAI|�;�����*�b�x�ء�1PF��(�)������.eT���b�7��>�D�����Ƶ�F�j�C<���|�A��ЋG[���.���Wk���}lk8>l}���T�M�`-;m�<�r�b�S�����5x⼤ZvB��Nc��Q+����!�tf�M�[:�P9�?���<֖�4n��GTC�
*)'�V~��·���˛�~n �d�����M���zw�ˊ�����Wx|*���|�����de�Y�F��'i�L�x���T���+2�vV�G�E��ǖ\DJ��2iJ)ڼ����$Y��5������km}�&�N1�!��A�>\��`�%�a���ϋk}Sܯ�i�z$(�M��T�~?]�.�/'��w��i+�I��lX�{&p����!H�����z  ����I�!�gO�� ڗrf��.�Fbb���25k��z�0�i�ǧy���|� ̏N�Y��-�~C҄~~6i�Ï6y֧������`�&��媜�l�cl�qq"�Z���*`�����b���;�[_����
���Z�ܩ�>��Jp.H�]d/���bidU��*�R�D%�#H�/K	R�]j��&�:C�<c�ז�<�Q����WC�%�>��=��p�v!�U<������Xc�)�u���}K������E_W��kMX�O��@���Xz8���ݷqC]5U�1�'�?#Vj�=r)Kv��^ؿ	��U�2_8����q�*x9����$]�����1-.???��"CF�z��/�ԓ�Zj5|mc�k���K(�i-c7�BHk�Go=_��1�#��l(����WgKrRt��yܖ1ĭ�=��`���\��oCN�i����9��޹��1\y���!M�,���W�\����9Ϋ��:��G��W �
�e�#_���e6"�."�f�msl�q2L/2e����я�櫻�]-ӛ��6��ʜʽ����ivA�W��	6x9����	0�SBT�b��?zY�e��v����g�&o�g�	�D+62yg½&o���X�*�!꓈��Xt��{��4�b��z�jgE��>JcV X�PM _f� k-�7$��<�`#����!k\χ��׏�t�	=W���+c���m��5�~��^t?ᎄE�S�2o��{��W?�$vy���&|�Jz���q�����f�r��en�=p����l[!����� �~�([���lNH���;ƚ�Xޘ���5E�4�}�8UQ��C_��(u�>�S,7��-1�-6Z�������1�+�Kb�@�<��XU! ��r�#/хfN�d��r��݄�C5�3:tO|�tx�eSE1�vk0 �<�0���MO1�j0�_:�ERJ�h0�6d��z(����1���,`�P�s?U�Թ�a$ڤ�����WK����J�}��`l�U��+��3�,Y���]���0~�����i��v�4B��`�@�x�!E/#	��]ݣ#�-Col���1!O�}0_�E�wj�~%�T� ���CA�#y�ۺY������x`��u=P�����Y����'
���I?��5�@����k��	J���u��x��;��}���KS�Xơ��=i��(@�Y�����T��N�+~\��qNd�o�%���n�P�s�&��hˁވ����r���gq��s,L{���2���1��cng��Hy~��~�z�w�q��1O0�J��i6��/�2�6V�����Z��ܢ3.5���KV4FcE	r�����l�y94�Ë�ѢY�l�#͞�S�J��}���1B��aF�"~�`�w��?4�y�%s�� ��G�&
Wq$u�Z�.��W�ãa_�>}�e������5oC�4��*�Pb�s�	�����]-����x�BN���MX9�ؗ�8oB��n�����'�����N��[UC�z����*Sx��fs�-���UwwG�J$�u����&2�Q��"��3��p�x�T��c�+�7�����v99
�W����A��λARx�_��~"A�_�!D�|����ɣ���<$��2`肗p8��u�t�ElvJY�\���:�5rM�Q��Φ�7����2����o�׳�-�A�E�D���8��D��HX�R�b��7D�L��I�!������@BB��J��K�y�|��P��M����W�mz��S�F8��{V�i<tb羮�Z�Ǳ�"���IY�p���Gp�0�E�x����q$����|�TK醊���0������E�~D9���I ��EZTO�����p�-`�E�N`�+����h�3]�*���en�򛎌�`���<+�CR#������S:��L�y��p����g��>��J��C3@0�F�_l�C�Gͥ*ƴ��f��F𞁍vVVV��s�p�^qh)���6��vz��[����t8j#�����RN��Wu9�nݝJ\���_�'�H%/4.e���J�Z�Dc�~r�y��Z��	�����0�LΘ�$���Ws�l�e<�;���5Rٺ�Oн�R�j��g�T%_s{ ŀ�o"�m+���7�mށ��*T��-n<��=A����ϫν����.�d�!r����mU,����������5n��o[%Z �`�XiTDv�A��$�ˎN�s�lw�n��#3Nf>MY����E�� ;`	u�2ľ��:?6-�2p�LʮS�{�����`Z�s���X��M
=�:��c]Q�Wwu!y�+;���Eqb����)�m�S�}�:���Cu Q �/��RX~��:h��TePXQ	�y�w-�)Ti�s�7YM�����g�Cc�dHkwDjȾ��~�>zA���@����Ј}�A"���ţ�+�se�딧�,��"�ݏ�����~^		>QLo@�X1�*�<@����}`r������==e��~��g���Zfp�����TV��Qm`��.|�w�}���LZ�(	�͜��<;�m�V�	��+;��2�N�B�EwW=��d�f��L���I��O!0�ь5�6�,� &��v�̫T�d([ ��� ��\��D�#kG�g㭕����OK����he�*�RHo��2J�\�N:֫���d=�f�
άN�D9�e���U���]ߍ��j �%�I7����a� ]�E�c�@0r��Nv�>�����-��d����}��Av�<9��fyt�^�����[ndl���5bb\8
9�-PH�*0.� ��S�>�F�ՖT�h�C{���B����.}NI)�"{�,�rZ�R�}S��-�Oo~�B��z���n������#o��Wu���� ��5s�
ب�t���~���6�$�Z�ݾ���g�GG��4|t��OUl�&�p�/��M�ZOQ�^�&7ܚB�R�������ʑ�O�6�jAz�����ŧ����9+�7�t�N�צ��RǇ�?o<�`G�W�ӿ�׋�,�s�4l�9A; �3]U�Y�]��~��#��
��ԑ���c:��,e������L	6^fR������G�g�)
ea���7�'�O�5�*��S�ͱ���K��u��S�b�e�-aj��E
�>� �fX1�V�qà>N���:���+����uv`.1i̷׀��;��U�}�3C���en�U&z�\3i�I����y��z�T	�Ǝ���rt,�u��r$����N�,ʟ۾<B�"',�V���Ӈi��V�M]$5����D�QLYW�(�����뫙��'+6����lx�4�m��TF�����)�9�3�1!�S��_O2J��U�l��rO��X��?7�6n��a����BH�6����"D��o�1�b6���s�b�������n/E*��M���u
��擹��<��E��܁>�=�=ʨG)��IU�,MP��
��%�&��/�U��=��C��<�JȻj'����]=c�pA�C��o����|/DLP�Ւ�o򠭮���?W�
�A0�X_E�<$�f/���^��ZIɳ7���Rdq��+�	�Y��KҰ�@�Q%�Q�l��g�F]�o���7��Hֶ���E\�P�m�Ž��������۟�74���o�����(t{s��@-��l�v*����B�ANkk�Pb%�����g~{؟�8�צ��'�7���;W����I��	\����q���e
C�Mq���,��d��,���^�4��[sl��6U��Z�F}E�[�G�Ʒ���T��A0K��؊��]v���}�*x����Q���'Q��%��9��an�`�W��ϡ�7�K��\�_�gTBP5�\u#���y��K]�C�.��f7���_��hX��	˧�2LT�H�ѩjE���S<q�L�:H�H+�N��M%B~@�٧c^煈@�
�M�U��3�?���P �d]|�n��]f�L���8C���-���e�g���F~@,~��]��MY<N���ݣ�K���OO*�Ѧ�m��K�{�b��>���T�{�iX�<�z��� ���]��d�6�֘�X� �U��jX��b�-��=ƭ���Aފ�����Ԍ[lz#:�s�������k/�υ�:�v���Ƀ�6�48N��1���+Y� ��X�dx���L�m�at4_6��sǦ��64����oS�OӼ��d��S�<�F	����т:������{jع\�w]��`���ߩ�C��8:��qw|[���J�[��E�F[J;�m�m�0p�6�ĥՒ)�Zi�}�f)t�:y'�H5m���AP=��Ll�ː2���h!�-��
�2��ϱ�!��t[�\�u��|�{JB�
��{Rv^���;?�(�mY�L�]V�rE`�#$8$�b�	�b�t����q�"&���&���	�6Ӯ������*�U�<����Yn�9�$�Bp�^���f��
^��nFC�:h}��/4�������ٽ�n�y���fQ�ʍ�zJ3i�L-o���oG\��U��8񎴉�����n��UR����|}�p���"�J��-�U� ��O�K�~���:������� �P��g�'){�����j:>=�(J�.�$�Y�D�����cX��P&�j�.��0��^�'.�@��$��O��vĐ���������4y��իtE~�c�P�4�֑���96F������!����k�;���S]�>�����'Àh���N��Ø�5��ힴ���c�B�@����3+
�D�#��	u��K���fLb�~ё󹕒����J�ρe�U�
�O�M�b���?Aߛ�=Io�����D�j
��UR�Ri�U b�Sġ�5i��^�)�6��$���-����y�bj,�jip�j�-��TEx�t�2^�<�[�Qc�Z��g��x.E�k�<�U�%���j�Qg-�3���TrvF����n�G}�111��ӶiB|�m¢�Ƶe�<𺜼H�.���_-�a�f��RuC�Z�B\$le��C.D�N̊�9HzطL�{1 �30��7�� 7�}3�(#A�����[�<�bЦ�QC���zz��*���g���(J����m���v^�?�
�eq��ӫ{��O���9�H������с,��{��&�g[��Cq��{�ovj�ߘ�gjz��/?��~�S:ㄹZ��_O�1���10o��1@$Ոl����Z��I�JM�=5�h?�lIoR�F��Z��ma�%�A��v�.N��Q+**
��O��OLp��y7�hcj��Y�Q���v�<���=�!� ��͋E�k�iؓ�N������?-'�9_~��^�,�cvr�#�,V��IM)��D2[����w$I!tr^?1?O�b��*�3��0��g׹<�>�y��}-m;1x�r\ �I��f�c��z���e��%�J�����}� �'��X	���}pe�_e��^Ϛ�i�6��V5�~�Ү����}����t�>��aBA�:Gv���@.l30l]�~]��BeW\x�[���t���m�������CԮ��B<*&�E_x��J��J�)���7+JUn���$�Q�U��_�6����5m��l$9�s���PN�  �>�:�h�[�ҵ�>��.��h������)!")�ە�Ʌj�Źِ
¤�&���P��=UD��a͐km���K�Ab{�Ql4�؜�ڃD�-:[���-NY�4C��M��p���!]g]9fPH/��̨֨�Vh[�N�aW5+E� #�������q������2[��w\�A�V����N�Z��k����v�R���4��Ig�/?lW_�;ǉҔu�7
؁,GU��e���j�S�M"��qr$ !!Y��\��b0�-�r!���'ӫA��n��ޣ�*�M�o"C{"��Xh���T7�u6n젠]�4�L����\H�ږ�����$����}P\Y�vXoSWz'���a�b��l��a���+6�;����87e9Rt5NW��K�aR4�?��3|��p�����z/!�T!&V?q�UJQ�����l�[�\�;Sns�֏�M^������|I���Vةh��B��cծ�r��J�`���M���Ɉ̞�o6�������{`�F ��ΧI*@ ������B��lw���?)����wf��۞�*잕7,��T�6�)�98���������
����nO�x�S�����[�-��)��� 3p�6)��`ɀj�үf�`"I�A�g��H�Rg����#f&�t��O��Z�|RD�e�1�V:���v��q�S&�0oQ�+�ϧ���;��3�CTҐ�ta Kvv���*|��[��(��=+�����L�ǤA�n�xUը��
��RY�����	�q��Q-�e%�	�d�9꽟G��1,"G�Ć4��#�F�0ө=O�jVW�>F[F8�'�c��@��&�����1}t�� \-��am��;�����w�
���:�d,�#u��¹��L��*Vw?���0�78Zw����o?�����/�e=�{؝���� ��������W���
3,IќM���y�Ly�~�=qJJ�YV�v�C(M�XJ<5d��f2^���sv#]S�8� 3��E3�N�J���t��g�v�N�Ce�H�/�J� ��<�]�a���2�8sC:�*''�1�˯"���QY:�xha�/Yt�Z{���Z�"6$b�X6�~Ř։�?R�����:�����7��W
Ik�Ȍb�D�6�tx�{G��e~��4)z�5�um��^�B�߅w�.�_%�֖|
��Ådo*��-y�q�F���Ep�}��߄�q0C���k���!x�NB�ᦊ/d���أ�����>!t{k��2f�QH:aD
��-�k�q,Lo��L�]����S)#��� ��ڃ535����q���0�3O�å�mB��˘�m^.���.��q�g(o�a�.���Vu01���y����_����f ˩*���珕KR� �9ϯ� _s�n��<:�=�{�ܥ���Gß�P��<[�i���ޘ��r�{��2���9��Z8NU&�dF.���R�DE!z�/Z�ք��L(�xY�7��;���Eo: �&6�/-������=a^�r���.���m�F� ��C�b�b��c�%��i"_������]�1��*��<^�b}�K
,��?)�g �{O���=?]��c�"���,LLȠZ�r�p�h�b!��u����u`wG����R�����q��x�u�7��\�<�J�����'�
8���Sн=f�A�9>�X�l֧���X7x6:/u�u9��Z}k,Hi������G�����#�W�~zF�����iXbZ\oxg�k��N;�6�ھ���ǭ�큦_̙�u���-�;>>>��Yh� �V�]quqrl��_ڢgb��'��K�0��~��ȇ��Z�:�(�(:]����0���^�4sR"nޡ�����,뮫..��.>B/o	��jN����4����9|31}L�4u�����q_��k�:����:�6]�L�m�놛6��~�fF��j��M�ݵ�^n167���h�M�� �~�fV0��T���h��t$��7SVV���{Ubw� �z�"�^+қ�L��77���AtT��<N��p����y��ܮM�pŅP��Y�,�(�Lh9�A�Y1��;�H����2�M������/.T.n�m0yѼ_~�皎���o�p.3m_�U���s2�W���ڙ�s�u�	/�˜D5|�h�~��~�w�2�ˋ3�����l"[x]I�������k�o�q��̓'�d�ٹ���)�\���f�\�+��0Y���y���c������;&(	cWg2pFmP[_��X����N.�?ɣ#��!��:̱U]%q�YV�&���3h#A�9 �K��lx�
�|�:9����j
��ƒ����/���1e�J)��,|!���c)7B���.�OL�Ȁ�e'�1���n]���퉭W�xǩ��ô����KF����nN����������P���;�������x��KtH&?�~��ch��K��n��^f�6+f��`�2�K����0֥+Y�$R#�(I�����y�~�FЖ�!ßC���X���_�_��A�Z�C.�$zFn���HJ:"�fz�G��*<�2Š#�g�.���&�%�)<��sC���qˍ���d[fB����n��~�������?�)6���I���b1���j�gi�o�����	�ra��j�&+�m�n毹xe���d!��Z���D���Z���3�l*�3�gߐI��>!'�E�����> ����sW�Dz�w*&���p�(�T�#	��DX�߿Y�{2�\"&�<g���D���l�?��jBKA����w��W�)����o�R7V�7���Gc�u���¾�4l8�W)�w#��P�����
�ց��ų����c�l�^s���虏���H-n˖�L�P�� q�\Dv�x�^dٍ����|�L���e-<�p�[�+9�����)w;�S��N�E�%���P�{}R8�@χP�]:�B�v�V�7��W����$��he��K��e"����LLړ7^ͼ�ط�C�|�u�zy���chíR����r�i%N���!��i��5��&���vgmKp�	��H;��hgwsrח��jM/D.�_^J��Kb��ElP0|�j�$b��wfz��ٴ�zn������p*R��?��2.h�ͭ�{
Q�^�6o�M�����D�!��ǀ07������cg4�t'���:���j�$�,��pdaX�\<:��a�G�1tod�i��9�:�w�]�M�u �e5��+�f�|��e$8�H�ի�и��{��vw��b�+tJ�x��MV#��Dcd�V6
fR5�@ �Σ���p�Ja1K�@��G�s	W�}���x}�����!���C�6�u������/�σ?a{b�Þ�_sZӿ�Z���}�,�yu����\ٛ)%Ƀ��k�U���)V�k�\��<����y�����u��oˁ�1��y�e"��✆?���~e�I>�r��_���#�������O�?�l�Q)��'�vk^�H�;�dgn�Ъ�����VV]���+jj·,���M�H*T���H4@��*�kMK�̶z9��2�\���rcF+�4m$.|W�ɋ)��bL�YGץ��l�؏�i%�?`o�B*��~zI5%|�xV�U��b�m�*���i�=i������v�����G�\�|[����d:.H�b�߷u#�������C�,іB�X@5� Zi�sX>���W�
K��8����.��D�G�ə��l�*�k�#��90������,� t�y�*;:�h��=�X���G��xl��W��_c���3�y/�;�^TH>�x����O5��PPPx�X���TK����9��<D����.�%y}�r����#W�{���l���7�W���D�J�9��q���2���\� ח#h.�zN?��_�h!���Y�L�0$:z���?��u$�ˀ���M��HL����7�㈲-�C��i�8���p�����⥬�L~Fm���f������?�t���Ny�}�F���B����AkB����/���G�Cm-K���m:��: ��7�[~�/�}^N�o6�ǖgM�=��8���37�سL��Y���G����]%l��"V�b�1C�����r#����-���#!��u��`E|f����W]3KM���������(�i���V�Ux%��:�����%�=+_�����6�p9�0 �~�~-e��Ʈ0}�9U�w����@�
ם��0�eۓM�雚|���̻�r/WǮQ�+���6�����˟^�0<�II|o��$�T�j�:H1�g�s������7�����Sk`NP��Ş"��0�O񴿶�Ɯ3��[%vbJ{��K|H�����T���=A0wؚX\n�H�B�׿:L����м� �)}0YD� ��J�+K�Y|E%4,5�]7KL0�t�uT������V�nI��a�������h$H�4�s�HJ�V@R�H7�n�����8���w�wl;���}�v��ڹ���֎ϝ���s��H�p
�1�+)X�7Í��kIN�7��nb�/��/q��x��"����c=�o+7б�8��3��p�%��\&��}�-�V�1r�TH���~�[O/r�\��}Ȩ���z�{�-�Ne�/�I�_hk,f���`��L�I�\B�zmؕ��`z���1
i�ٯmO���(6>^,δ�m��k�3��½g�MMr	�X<SJ��f�-c]Jܴ��%�A'��	��Fe�t�n=�T�/���yW ^,j;3�6�J��V�?�e����E,ݗ���Ð���ϓ�b�����;}�Y�l᠁љѐsa�H����Oћ�v����Y>P�������0����x����77��״��w�?3V�/���X��H�i���R���7��?[������i��ii��b1�8�"ù�X���/Cw������ՙ��h<��us�,�C^�F1�@</|�9]���!׮}2���dA��M���q��N<;�@7�rէ �n	7k�ԓ߁�) 8�WαW��Z�X�E��]X����F�@�Ȅ4%�Ϲ/2H��Z����}��]��{�%_M������������
y���:�|����hn V�sw%���e4ِ�ce8�qbxD��ߜ��[N��}�@9Lt�[�Xm����Q��`iF�r�7`h�����@����h�`����02J��N��[ô���;Tц�� �T������X��m4���T[�ͱ8i��1�(E��(��\'�=_���F4����\�d��꺺w�7}�'���ق��G_n������E�t�K*D�q�ȤY�9�zcu��� �g�dy�_d<N��Pk ��{���3-��[�̼�g+#҇"mr�F�$��ۂ��hb	�jB�c��/?m�]��7��|g%N[�:L��J z5Гw �E7��'�>x�g� ��益��ZB�P2%*�b�K^1�"�[]�=���U��N.Ԩ`���χ�8:�wD ��}X\~�(U��b��M��y//����?�w������j,焇?���͎q�]/�������4��6�$J<Y﫽%��8��2דO+��=�
�4���G��w�YW�RƮ0��&����A��qs?9,��қ0��j�F�g�#�ǹ���n&��'i�+_��Ɨ;�{����7��%���YF���݁OlLz��/,�屑S���R�>oүLf����u/�����i,��^�	@��%�<�5`2>��+X��8��<A�Ն�~!�A�sOR����B�x����j���$��:P�p�n����y�e%p4D
�_���[&uap�D0�:�W ���}QXɇ;�ߋiӮ��!�I��Iƾ� �����_��M�/�K"����1��.KF�83s����fD�~�J)�,�CٹY��q��.]���V�5������5��e���wF����
��D:��آ5�gd�5|����aO�{	�[>�GR
�a�����d��j�ý�<<¢�*��L f�U(>��z	��ך)�-�r �^�z�*��z6E�n֪Vm=����MԆ��	t
��5��n���xK��@�v�l��h2�1��f&|�p>7,S�~ ��Y������qe��nX�.F8��Yj���c�ʪ)S�-8X�a���R�qh�����w7���h�)\Zo(�p!%������-�[����%� e��jF�Й���p��p�uA�]�����,�.w<�N��a�$N�Vk���,S��"U�hըuo�R߬���O߳I÷i��R�����*3��� Ha��ڻ��=CP�"��\DA�.�*�i��i���"�3�q�t�F��?��Ouda��XZBI$�,�hH�C��1�n��*������R�`����i�:������%N�Kt��i@h��z՟�Y�+�@�i�m���Q��c��n�U��uL~��L�a���g�w@U���]��C7V���k� ���^��'!�4xX�?z�㶗�q�*nX<Z����z2�X3;��Ԩ��zs㎞jd����*��$`fz��A��z�N�U����Nɴl�![4Ӳ�����"���G�=@=�&�S�S�h��ui9�L�Zz���9�Z��l���pD�����K�I��|����e_�BHڗ��9���v �Fq\�;������ILi����7�נ
��nbR)J���������i�e ��0U�UӦ�z�E �r�O��7��^:��J��TF�w��M�:I���ãa�Ѫ�x���ґuR~{Tf$��/�ʋ� �ejL�����<�߃lٔ�3\Rƣ�>�_�⒦U���2��
��r�@�ܒ7���32�M�M��"�]! ��٘������܍ �_Get<_������Ρ�X3�3������t\zL��~�zF_zܼ��Ґ	�\FF��Eq�_�~$��E��'i�yLhu�>9u��S ��f�y�y3U� ���[�{���8���%>�W��L��֗g��8���3��iVv��0ݴ ��C�O6/�'�g�>-S�3H�����Acb��=�\����;�=B�����ج���ƭxm�X�!��e�YE4���1Ϩ��P!uC�̌:^,������ ��OL:c/>�Ĺ���%�e� ��rШV��m^xx�0P��#����N���]%�7@���Y˷|9>��'s����rNÎsM��liGR����Z�Y���_S�����B\������_�o�[����-�N�ژ2�c\>��(4���u���sK����veL��A5ټ]G�wUi�ƞ:ug�U�q4Y��8������3�T�;m����"w�&�bM{Ҙy4�����9+0�W���n�֓�v�g�ؚr�Hı�K�YH4:��\U�t���q��H-r#%��|kY�s��$�N\<�g9�Mwn���x�tS�x�/�����q�\S��T�Bu5׾i�����6�na#�J ��q�I�o�!�<�źۥ�[����ʱ"����ۊ�8H-N�*+�J==�G��0!ڬaU6���F�A_ק�No-p�.���p.�!^i���q4��8�	[�%��v�,���H�z簶�E)B��/X�����w�ia2�w�.���X���������1�faj��΂��-�Y%���}�⁨WV�.)>�+my��+C�i��Ǻ�o`��@g7{4cත��P=��5�e7U�u��{M��u��XgZ�Т��(��N��A\*��� Y=�-��m,�0��4_8�F#��6I2��q�$�$W�\�	�T$gɸ����}e:� Ey�*5���h��g���aY䦙�DJ����3-@��'_R�4M�Þ[I��"�G$��ߒų����L�wc�"a����5�G��<����܅���_��wAy󡭑'R���^s!4�\��j������;k3����U�0�,2��s��z/:��o���a�X���L�R����&���3qL4�j�0�H���طo�4��P�h��z- �iL:��鵌�s�O	�7u�YƠU�ove�������i?a��O��o��n�����o���)Y���I#��P����${��xG��q��$�a�Ռ?����{�G���4B��1m��`����jg^�+)$��8�/��rI���B-Teo��r�m[��*#��gp�< �E�PW��e�%�^ɯ�z� �akƃ0�gl��Y&���vf��%j% �x���LA�~]�yd3%���L!SS�I��B5�N�ϘO�XYř^��o|�GRD�c��)�����E�/*r1^�!t�;njV�L��J�hf�}[��g�L���>K`�.t�A[�Q5#����ˇP͆���m�$vV>!��H7p杖�~��*�7�
p���~|7�9�$<z,���=0{zȍ0ԁ�cR���WyP�/��0���؊t9�r�$�?.[�~�wl�ʢ�BX�]E,]*�G��c���t��(`�`#�e���2� 牿R�*~��pj��֢�&��������n��``6�6�Z��T蛝�+!čRE�	߱����[7�޵e>"h�&�;���E���r�E(٠L	i��2���L�����4c`F2[b/�x�4�|B��T;!7�����`��sJ��/������'����c�|��T��e�҆���zx������lPl$O���)b�d�(��
��H��9;e�*5�DkqN2��40DmV�04+�o\��6s�������6�`ߋ���w����90����ʷ����U����jBDI�|��N�K�@^b����;0���ƋF�@�~q��#�4�a�87�|����g-��M���,1~�/�ڱ3B���x[��Xv*��@�R����s�*6��Ջ�d��>�A�$ ��'�w����%�0F�hJ�1�L}//�ޑ�~"ヸ�>��i�7&<��`���8�%���%�"M�H��D�̈́�O���i�0W��D@���3/�a9�d2���)�d�����W+>�eHN`�I�"�w �@���W��	7b,8��rm��1���P5������Å����zkB��VJi46�*�S��n��w5�o�Gl�l_lPsh�� �|gA� ��G6�O�����MG�<ϼ/�*��A�p;/j�L�\��$��}mD�89��_&��0c�w�9��Ǿ<1���<9�kZ�_1��1Z�9Z��&=J�8vI�>=���^!��x�ҩ�
���(0D��R�b�#l����+��՛����B� "6J�X$Z�87T��7�8ǀ�l
�H�u�K8������*|�b���[,�<�Cf� %�Jo�����x��s�b�����G�PX5�yW�����.�"��*e�Z��g�ƍ����)� 5ko����D��Z�EU��Y.*�p��RMz�@[��vF��s��QRy\�A6����>M**��)[�����P�.�>Ը�Z�74�k̄F��Ǘ.:��nM9հ�n�h�����݈���H.�16��Y�ćhuO�ϙDv�f[��$��W��,J�A�C_��_���G�@��3��/���ئ�us��2��|q此؝�E�f��������PrJdpk�~+n�<���J4��4�Xt���"X1"eMF�O���~@����۶�0�ף�G-�?c3#��3��6m���eor���C����ޏ��S3e�
�҇�^p�R��=��7m'���{p�E��;Ǳ�[�?���z���Ur���u���s</⋇�kp4ѣ�r>�J�sx�;��g]��ж\Ȩ|�'2[�����ִ�o��a�!�V��{.�G�
m�<����L��ih�ϩI���JR
x�iL0�g��ɴ(M�Q"�`}�PY�s��ֵ?�1��m�{��ҟ��PVgS�Ow��bĩ�z�X�+��[w���^8g6K��"�ƿ��y�FG�z���y@�KFx8]����%12��y��z�m���\��n��́����g[�&�f���x�cS�����MOX�~����̃.�5��Bt˝I#��>6�7ӛj�] [��;bv/_]�k�B���;XLq]VZ�:;���:rP�v����/9l��؃�<fi�_���>�7,���4����h]d��p�m�,F�:$y-�t�Zy�:��g�{Pg�=ɥ���ۨ&@v:�P�iۡ����u����T�;�&��?��A�=�J�6(�����b�����ޯyK����jn$��v��J����Ss��QEm��k��xT�"��d�M.Ǵ�����tv��Q�rd�����@'6�l�V1���u��ݴ�2/a+]q�>к=`V3*����ឭ+wk+j��bu��aJ��Rt9�j���$���s���g�TO��Pfx�z3eN%f�ݘ�r��[�jc.ܵv�C���!��k�UKϛ����sS#��Z��8��M�<y�Q�r��X+\2���g	z�o
>�bc�_�)Rg�T��x���S���{Qd2�;�४}h��4�N�<�ʨ)q7�
4G(�@\+�.XЯ�)� /�:�ZRN"Qt����ٽb�(d�E���q���X���b]S���3n���S�§��㉡6���Q�J�ڒ�Y{57�Eu*�?�ֿ=�o�����s cy[oզL������n�sT��l�|uĕ�g\���Ý�����ݼu����'������s�@�yL!�������;��=��z�G��o�W��8&�XFD<�&��l�<���Ӯv8zۼk��?��ϝ ua2��[k�t	 į�ܿ��S>��j�Lm�����z�y�GgY�,�U�F;�f��RN?�샄�m^�j�H4DW*03���%~���Z]�.���-X�%F�2��,�8���"��p�p�ˏ~�xP�f+K��˖+��a��^}է*j�<����j#�=��������p�����	���s�-�/4����"�#וʙ���:@2�M:��DX�Yk����m�6��ή�g`n�Iω�zz�]s�{h��X:Ţjo9�.M8�"���yxy�����F�:�ǷÃ��f�|?_Ќ���l����q��cȓ�hb]/y�#��"�0��a*�����z���V�,�o�~�QJ������^����cF�m,P�D�{�OV�۝G��r�;��b:��^��?9�h�"�/�4���Vl����,2}�ݡº|kq�1���یA�j�2��+���� �*�ѹ?i*5ڝ�d�I2#If�z�(�G|tY����-G��Ig5��ß���?��|&�*�fG+,�3e�?��l��&cB��΃ݚ���j��7�Hֳ�!*�}���\����R���-u�߄$��|��&XS$JV|^�%��B4��f06�c�ڏ���,'�����sH�g˚9;_�5rH "���X�����?���+
��&�QJin� [W���K�6�S�	i,�wJ1��ֵ���-��c�_
�>��ǋǡ��[=��YxDm��F;�[U��4����� �ڧu��]���RР�@��x��m@�3�i%��DѾ~�S~jq{�k��㧀_1��p��X���csإ`�O��xy�&zt<>k*E�7��3�|�o!-�l��:'�$FMΚf�#�1G�uf�<��0�K1��pb�>�q!�[]n|;�\��~vN�K_�>��꫍��xj}>�RچZЯ[qW>�b�D����V�[�2�ݑ�������1σ3!r�}��'m����/����&ݿ�N�A�_����um���.�S^n�r�jq�bB*a�V�S��
��rG:�"��"���cً�g�L)�I<�+�ܹ�?d �c�ؑYO�V�|�j�B�o�א��
i���S�{���|][ޓ��/�*���H�S�>��M�[����K���a�ߝ�m3�W}�85.
�>aHD����KM#��1�:��#�Ye^"��/^SI>���XX8����4�����Rb'��	���e��CK	w�Ec�ּY{�͇�)������<�٧��q�a���C_��4Խ��h����bZg�:�"�z%�i�����{����ͨ�F�|b�K��er�?�r4U���I�T)b�N�1�O�<��qn������{�p�b�{��d��Bq���V�;G|4��t�[��B�r���&x�p?y����i��n��)W]���6��&ѧ(��"�<Nlh������8��G�#-��h�s k1�����7#n�k�4ԓu�!РBh~Y?k{�2� ߉�@d��&3�,l�H�J>~�ԸH�W��1�KG����ȘayD6�2?�W����?(�̫ǚ���im��3���D:�˿*��)f�2��\Fҽ]"7�6��+QG���9�o�2R�Jg�3����Y�̄~b���~Fˣk$lM����7����8����CȊ��s�e,�|�=�^R�f�m��p��y��([p7?�a�k`��Y_��3��>�ZN�s��=G�R��߮A��9|e����~�V�ɏC�H�r�Eg(x�����V�1�3S�:�#ԇ�%�4r�j���@(��?��y)�KCnF���a ���J-GP�x�M��tQ�e�'&O��uz�wT�HXσe�$�
��D���~Y�;��\��M:|.዗���<l?�����*�\���᳝���|�K�jI�D&�+¹�������
������y� "J��)f�_(ih�7x4�N
��_�o�7ڦ�i�f��_;ڑ��0�aCU�� BtT���(�<�2v����Fq>\�m��'x\@V�x����9�%�S30	�Ufm8������l��o�L�,�4]�k��Y�Kf�f���/�eŃ:�U7:K��bRM�$���/X��*�3��
�ޡ_�=�r����,�3�L�k�w
�,���4wt.�\�e����9�K���Tp��i�ʫ�ܷT@���P���|�y�	f�D�fN�#�����G9��h���Kl;����*��7��Fb��=w�6�>D���`"#3k�*�"�x�fV&oF�6v(v�&&\=���m���� ���Lx!R�k�s�.�*T(�W3F������i$�ƃY�
o�%6�<�Q��0�y�1����=B9��@�KJ�;cT��Ǎ�	���mk�'S7W���|�	���?��qF-/KQ���Wǰ�ę�%������f�#*�Ԫ��7�o��Hn_{�U-l9��PP~���B�ԫ�ț,� �:�] p���d%6q̊�r7�����͆��%I�:��&s�v��_m���k��y�Yo��E],���	����u�_z�8��u���%3��k���թ� L��ޜ�g�-#����qJ7[��G�꤬[�
�.�1A��"��@0;�1+/d�Q���249��)���Xs�P#$�t��47�6����M��l�� ���C�����kAw3���3��jIUK��x~���I.�Q6�k�,��4ph� �zئ,	�L8�y+�4�G��H��6��� ��l��O0�ٷ��Bj\2|�����a���Q7T��f|��S���6������.W߂Q��5�P�e�;ϋ�����I员tby�sm�1E����=��+�k���"�f{s)g��h���bS}�`�'9��xq�/���M�-&i{�R�����"j�X9�!�\�d��k����Σ[���d��P|�J�/���F*<�!�ō5Ю��"�"���U4��-O=�<{��,0��h�u��	\�����D�;�T`�NP*2��X���k����f>�LZ�#�����:��`�(xϥ�0 �0jO�pX�s���*�lO|�	�xu�X�޺S��}�B �q��p��?3���=�_�WVB�$l������&'K�+d�qS�߿�mv���s�cT��uuA��)y�"!DYFcFy�ů*bΡ�o��:�o�ig3�Y>�Ҏg	un�}s����3��Ag>�R<㘊�Q���P�����ՈwCS�"��9��;U�}_��"��j���]������k�o@�&�U���*�l1>��6��s�#cn��l����3��z��|�F��ݘW����ʳ~-.���Ȋ5 M����G�LO�R�f��p�a��	a`�H8�	����rJ��f��Y���S�-��H�i��� �:S��G7u��u\5]?��[�n0�9c*,�S��$ݽ:�	����c�V���2������%jJ?(�+9��k�o�I� j���F�kH�*���Yy2ɍ���A�F�F����n>j(���矴}	I^�����\�?���D�U��	\�|��$��S���b�����w��u�2�#lt�ώHo*0{��;ku�2�}:B�ݖ�2��`��PV�n[hښ��-�����J'{k�!�R˰��t���C��d�ڛocj����t���%���j�D�&6\+0�w�2G7��R���T.�os+鬹H�l���+���ur|���Er��l�!�$����T��s	{����@>!~p���T`%2�3�h�JϓsS����l'^c}+,��݌�P��S��@ъiM�`��s���$�5���k%Lw~MZ�Y�U��y�Z�
ފ@�Gd�n0���bǸ\[3<9��ШC�QR%��۲{ԺI�P}L.g�͖��w0���<������
F,*�>S�I���dh�F��9��3z�����.�蛿XI{O^o��2UQ<�H�'SbudD맧�MՆ�f2Ƴ{=�/�'��L���U'��'�xf=S����i�5��o�I/�6ӭ��8|���:GJ����ot��ɝŠz`�Q3fBK�*:]��A��/:8_/w�0�R�rx��q��K:K�vH)
Bl�L��w��v:FJz�xv�:���ws '�q�	��;��Þ��.N��F��h��	�����>c�&�"4�s@�SYt�*	�ܚ#U����V�;[��?��m� ����ͯ�,TFM�4R�Jr���d9�H��?��~�5��Z��ٮ����q̬G:4<g�Ԛ~��W<`;������o\IH��������λ�q]vjZJWV-�����F.��tq��ÖA����x�z:����@�k��|*����v����:_��-��yr$9��K��?����s�z#�Q�`b��9^������C���Ӛ/n�"����5�Z�ڴ=1��m�jo�A�߆���Z�,��d�YdIТ^dQQ�1,+Q�̖9�ώ]\�K�+�j�@�1�<S���"o~t���ZY�#�A_�濅ͷE�R���LJ.ש�<�w��o�Mr�{a �7���\ƫS��&L��D������8�Z�%���V�*G����Uq�Wy�X^��&�o�ӿM�ڬV��Հ�<����rS��\ש����C�_~QL#ȕ`O(9e!vha�TK!C	�� �
O?B����Xq��W�@���B�}�����2�%1��2L��Y�������ɾ�&���:��2�r�;V�Û��V�� Ң4�P�,6 ��q�o�Y�4�Ŗ�!��}�d����P{�,]_��=D�<Y��D=*��j����iTcJcK�Y1��a�/�8���3+x��5�� �`bO��*#O�_Q�R��ѤFZ�����_d�]aC͢�EZ5��t��e�t�ݹ�hde���LV���q���	�m<��*8���f��1�G Mr2G��_�G�w9O���J�-}� S�'�A��O~���>�K"��E�����#k��.v�$K��9/f�0eq`�͇6��>�Bg�؍����=ZH+	8���5��G�P'�ąrc?��������,��H/u����Q�m8%>�.)�h�ʑ����C:[J\G�3��{��W�e�2e����>�o0��(Q�C܅Mܠ)��*�"&�n�������'���Z'v���_oo�^�a-*�f��>�D�-���a��%̸&���`l6��D7ŀ��u#;zՔ�3o��5 x-������{�J�I�����q@q��O@������`��
�0��p������G���/�Z_��8����$�:�h��	���+�����✟���}�8���5�A�E�w"ղ>�qT%b��t��T٭Wƈ���*i㈈ۈ࿨RU(>�C���� H���LX����6!���f<~�o?��>;��S -��	�������}�!�;}�D�N�l7������\��%"7�>F,�E>��I��J�97�!,u�U��S��ȓ�'��6���dY9�f��]���}�x��\5-��_%*���q��c:�-�p)���2⩙�}������x� :�Y�N�u�`2� D0�D�Y[����JPL��O�V��9���Qt��?�YN���?
��C�Ԫt ^�<'~���-2��1N�l�ӓ�Ҽ!�*#�DO�p�&�3��&����sP���H�7^:o��6��x!��,􄉡�Pa�f9^..��h�a��<N�^z�1��R��
��9k0���U��i+J�s�G"h@Eخ�|��HR���`�B�,�����G����N|?{�-�׆�j��c���O���:�����[`o�o}/r���*����Ql8U���h#�g�8Xߌ�_���Vy�н����7��9^�}�j����pf^��NGp��r{;/��BJ��M2WZ�!�/ͤ��~��dA�vvu#O����>bW�2���vJpߓ��q!RE��2�ߐ���9�=8���#PS�9���H���E��S�z��C�t�1G6��⤚��A�@{��j����x���܂W��o9M��n��]Z��!�o^e�O�Xٓ��Ak����u\�J�PU]�#�ͯ�Efx1��%��КT,O�U�'�V��7O��J_6*`S2���?%v��C��*hc*)����cha�KCu3�)A�8WN�����S���7rT�h����YTaز�x��7���/� ��S��\�i���-�^��/s�lx��u�ғ�BX
Nd�)��˘ki�>���
ժ�G('�J�u
��>O韦Gr�΢����i��-J��%�3M�A����^J.zq6H��#_��T%��*�r#&+L��@�����TĆ�O7�>PZ�`vD�U?� t��^�����R^ ���ĪｹϱL��R�.�@��2�'����܀��1������}����MCP���T���q�o;t�$�?�w<1*z'I��&�H�D����Sh�����dv"���я̞A^L4��vy�e"5Us�Yy_�<l�Z�ݻޯs�x�S��*z�����Q�8�/>�K�G���Ar�!�R��x(�2�{\�/�ߊ͓._hJ�n^+a�:/󐽘p�<g��o?����mZAGT	��_�Ӯ9�Pe)�05+�Q����T����!-L���
6�������: x��`�T&�� rf�)��Re�C_��YJ����^�+�?�!�r��z6�jJ/��T��P�7����	Q��}�vR��Ӻ��ةʣ�Z���g�}�)g�K\&��k`@0f�����'�7ώfGc'ofu����s�U�A�Q�\r�����8�*�������^�Ķ��fG�Z��	�Am{n��K�U3�����,>tK����%B��:[%p$m�I�����&������1�Z���obily�����ǪZ�D�  iGmԮ�����gH4�B0Ψy>OqU�*y:���5��j����b��خ������鿏��BK��G�%�1���,���/�u�`���T�L����m��Q�N��iiy9)k�/&��[&~L~Z�a�5ؔ9�侦�M�y������d�Ҫ|b.jj��N�W&eb�`���ao����7��l��ie	��J�@��?t� X}}
��`�����i�9R�)���4$�}D|<�n��x��c���K %N�;t�&�zL���	]o�����BZ�]YGfb��dH������x��˩	���L�Y��w�r�� T��=�I�v
�OF1��<T�}ИR�e5�c7]�g�k
;g�T`9O2W�]��0��3�+��(U�5K��cS��ӀO��K�j�y�5��w�+�dԪ��p?���,��1��>���7|�@�i��/��(�kQi
����W!��˄�eܠ��|~�gxO��4_$%�U�T�pka��w{����fE��X�A'�^ۇ�?�K�Д鎼�/%����v�$��U�ҫ5_��pl�=��A�������lX]vna��8D=�b�_W�x���g��Q-Ӧ��;�������ד�E����կ���>-]�£�M-�x��J]k���?��Ob&���гC�Z�t��zP�}}��e��CS%-�0Je|0�o�����5DU����)d�i0�Q�Qh�/�$�3�RĻ͚��]��R�Vy�ʺl�'P[H��/��-Ѽ<I�EM��&<n�B�|��D�HXgz�"�]�(g�O�	V"Z�>9��Q48��f~$��?���Xn Q0�]D��BW&��d�S����m�q񄣭����w�`(�X��>#��� �����&h�4��*�`S���UT��K��O��#Cj�ԟN����J���K��?�X�����&�MM�	���3^�'�
���#���j�<�{�充��ݟF��[�t��&�N6���ي��ϩ�M��S���|�镕,�Q��R�Ux��q���'+���Q4�E��h*BtcK�K�E�o���?��n��. �:Jb��?P��}��@LR�. ��$|ŗ]�d,��]���͸�s6/�q릎�����a��63��S)eϦ���p���B[�$�_e����3�\yY�� ������0���]X�� ��B3����EX�����Q�L	]�]yE:&&��Ƽ"E��F?�����Qt���|{l�#����75������?��쁀���S��Ge%T�"f�}�=���	�|nr��sݖ�?��A����;ܷ���_`�v�#��R��J���,fW�*婤hz��U�p��b5Ź0�q���{�))�D��!l��Ile(5��}����w[pl)��H�ϙ�,1e�O��li�}����ץVl:1^�6ԟ
Õ����h�a�t#���g�D�k�;�S��$=����A����a�!���X���!_#�ey�j�FarY1�A��\&������OeJ�Fus̼H���ߵ��b���Jf�wFş(�F�gJ��w �����ި��7m��k	�͵5�]ITÖ�1f�H)�8OV�7��7��;mu�}ڮ�{�����bZko8���Ȭ��Ojl�[�F��Q���,6��-n���3�ه[�m�~��h~��!߯?�jdH����� ��f����;./�+z\�y׈�M�_.��'�U�w� p����RպH9��H��}��el��8��CdzI����o����;�M�M��Xx{�$<(Ŝ�����w�b.��Na����&;]+�+�>
�PȮq��[Y�+�� ]����!�JQm����-RmRD��%��u��"J�.��Z����C@���q�wԗ����\鹤����� �=*_�z��C?�`z��k�N�i�9��|~0����uc[�hP@S��U�����������sb�Ҋ6��m񽞘�G����$�,��u��H&˵���s|��o�<�7�s����v�˿�&-�������okk#|���ʈ��K��L[f��y����*\Ҵ=?��9���gv9�;��nv�������b� �8�{�\��s�����Hz]^�|��
q*�`�SX�뙠X}T�����ud���&�2�p�9���V2T�wOr���.�M��X���[뼩�o.�רލAk���n��W�]�;��ws�7�>�9��<���vm'�[�+km���
�&%�΄�!X���)/x���l��$��]j����vv��*�f�8�DG��V�m;�w�s��	�x��V%	����;U�<r�L�P�O�`�m��r.g��5%Ĺv�wS���uJ�.EE0�!2���)�����#�Hӫ1yK�8s�FT�������w�O�:^/P{�g�}y�-ni���H��f�Iff (2J�c��t��Y�Yۜ���e&;g{C� �ӆ�9�Æ����O"�)���^�8C�_6;�
=�?A}�n>	�գ����T
�U��FZ�a�v;\pW�W#szƦ�Ty�L�f�:�߅���|��}Q����S} K(!j'�����n���%�${��~�B���c���Ov�y�QS���x5�P��ۿ��+�����$$�h'����(�Ӭn��?��h�9��d���̂�5��s4���\�8s�G2�&�k���5z��b]�������xEG���d$�B�e�@f��Je���"L�.A4{y�<���C.?��(�Wuo��-�X�V�����cU��	VP�3(*ի��w9�`I��y)[��J�\:�Mc��`<1�P��fVFe�~���7BӼ&b0��1[�9��,+a��]�L�`&�'t8w���զ�������N�؂�!vt��b��ozsA73ݛ��
��Z�NB�x�e����Ҹ��E�N�(s�kBPJ.�x���Iö�/<waXA�����T�G'�Θ6k���q������~<���<2��2���4H"WdJ<U��ڞ�S�[sd��>A�j����tU����.����kS���t��L�5�9��ܒ���i��6c1��Soe�u1�� �1-5���C)�t3tJ��ҍt	HIH( ��JwKw���~���4�ff����ڿsֺ��g�pڤ)W��}ͭj�}Ozp�����\��ݕ�_�[3����_�����X��l��#�R:��Cn��Z<yΔ��Qt�(^蜸Nd׌I/AM%\j�OY����郄�jy�7�a��U����
�.�I��O�
3RG>�X�Z��qe鏩�q��\!�����̤��L�����6�xШ�1���-1�A��g]G{"��3i$�]��O>�QY�oƓPP�Ox��K��e����$G��$T����{,�&
R9����m�����?�`s�`A��ʶ�/�L�l6���]C�B��k�n���w�քu^�u:�k*��K�'ɽ�����D��4tz����5~Y��I����>G_V��k5�t;X@���<���B��Q�Q�?��z��@d�w�B�3S�x�b㦗ZE��F��l2�7y'�U����/fa��=�L0b�OK�D;G���xvϻY�����߱�m��HڜhCY���_;�*π�4l����>�&�i%h����nt�>��!��Y)���9��/u�|OTK-B��98�����F_{��~����	��������°i�whҥ�H��(������F�h[��u���S����p3�"���5��q���l\��&U��T�[E�$J�)���ʃq�F�unC���BY�j�j��z�+�K��ꀐ\��6ըX��h~5���w���e�?��k�L5R�^�2�k%\������5D���Ʀ�{�ս	ro���fkҹ�Ʈ��嚵,CR�>����y��>ў�4�a#����=��"
�_w���T!�Q���1���#g�ں.�s�]�6�J�@t0\[g:<c�ÍzFT�l LW�����������r��X��93���&|+.��vx�C�L��I+�}�'����4U����Λ��.Ro��(��/�;��zU�w/��I)�ڶǿ���aH�+�c���U,�/t�pqgΩ�=pf��&�78ѓs�?���L~ȕe�r��*��~����o�⵲CcJ����9QR��U�_��&��� XjG�GB��n&dz4x�c͏V����d���;a�?��4�J��@�ʶ`�����Y��]ruD�T��x��tg�G�� ���I>V���|�$
�;���i__D�����+�A�[�:E��î=���7����_�+�<Ő�n!A�OZVB�=.�2X�컋�z�:	|�ȍP]q�.H�^�c���"q �].�Y"5�	�<��P|;���""W������mN}d��@�3��p
Au,�����c�� ������	��q��#���V��˦Ї�Ƅ|���Թ��C��p�P�EgՍ��2K�R-2J�5��\�8��oGg|˗���K+���;o||^3���3��d����6R���k�~]�)������G�=F��u�+�y�ܙ�C͝�}�$�|��pi�}n�ɹX>%�?X�α�0�`�|NH�/B���,��(��f���Ŵ_�&�k���N�Wm��^-0v��-=���X��5�i6>����M|Q��.� j;�I�O>@ ^폞xE�^2�������fݜ���l�s��e'�|屍&E;��{��ʃ��ud�(ݯb����j�����;׹�a, g��ʎ�swr�+���TX��G��S@/���fF�'w�E�	����P>�����'�-����	����9b2yLr����\�;��iE�t�����D�t

AP~g��	A�������4�����c�pRnx�\�\��2��q^�|�S���^b�Ɇ��4pk7�J/G�>�����ꦎ۬��k���z�m6�P�J��(��"����A����9�u;76�v�2W���;~�� E:HT�K�͔����l ��T�x�A���w�Ԙ��1��~;�'|�4�z^�]�d���8P�H��A�����$+��Y����"�fE�O#re�r��2Ḵ�M�v����/�l�W#�T�&m�������*)w���ٌ���c��Z�-*7�cB�/t�I0!�\���o�A�]0tE�-����#�o�\���=�9Ym��!z�t���3.�J���k�-ЈK�І��
�^~�R�&�H��1�$�751aɭ���<���j���Ȉ��y]+�͟"��Lt�>�*Z���}�jT��݀���;�q$�O$���|GS���+K2�~7K��X����R~^����>O>R������L��X{��'2pk 6"r���5|7W�j�(�����͖��Ot�5_r��`��x�'{↾N�j?tN��FХo�6����WfO>�ӿ�}��	������=�`�R��I�� ��%�Pe�eJ�'�57��Ju�K���8�;+?w�f�g�BcQs��O� z9�k�����܉�OV �§�E�V9~�B�!A֓�����/	��Z:����N�{"��w�Wʭ#��Mμm�ؓS���*������%ڏ��y��U��+;n��2����ܝm�L��Y�sy�+Uɋ�{vR.;-�u��;��qy��9�VL-��f�������>�lގl�'�y�XT��H8NFյ�O��|h�#�eɁ��6��mx0���q��[�����D��)��.3�Ul}k��Y�7�� �߷<5n���V0<g�`Z�g�� A��Y0��}r��1���&CV��_�tj06j�p�`���8��c����<��t�q˼�Ǉ�E[ۣ�2w��P(ؼ���nd��fD��o�;��1������* ��2��;�ue�d�-Id4�6E$���Z� �f��_ĺ���z���됃�f����d����9�Ɵ?�i�����D;����N��OR����:;'��=��1��2B���k�H2l{Xg[�����������./o�_��Q1>9h:��k����i �?����`+i͞�����$"}�^�\���Mx�P�U�ܸ���L�!��nH�� ��	zA��G^:��
gE�'g�[�{ӣ&�T�@8�1�hf4��*��o3}E��ګ���w�]��r��U����'U=�e뷽�YrFD&��)��\9�M��mofz�&;�ZG}oٖt�j�Y��-�����I�A?���K�
q)��@y��7<�͐���������L�D��x��>�]?��uZy���?R:6�Q��XF�1̵�A<��{� F4�������Kj�Г��}�ޛH`!%B�w�����$����w��~������b&<��]�E
-'}���A�z��g%��	�L��[�4�A���K�P�t���0�wx����Ӄ��I�!xw^�?(�X��\�ٹ��`��c���6l�ǝ0ٛ�ރ��o L��Y�hy��U�j��� ������v�$$'���߻i��W�\p\�zlZcs1�tB��@��z.j1l��g;*^�45Hi<\��2w�2�XC!����E��|�R����V���=&͏�q�/�vO���:��9F�h16G�`��Q!�7-}��9�;�ޟ�O/����2�	507��d�y���u��>�)5QfOhs���]�H�6{&�۷��{��&�.�9�e���/���B�64����������¥�tU���;5C��"�;k�T��ն�S��U�>�����Y��K9�e<#�I5��rs�!�8�D�+�3b&.�r񅋊�[�6[\��|���ih�y8�9�8uZ��_1��"����ƀ�6��/͵^�Q�0t��p`�E!J{��.Ry	�o��»R�3�*�5V��HD�����0'4��R�a�Z4�L���T���{s������W�yL�KWCF���y�̚�<���H����v&L��2�U����������P|G��f5VbA��G]3�|�Mi�V�$L!��>'��~ö�f#&o�����7G����K���������ڏ\�nJĶ��
x6ҮT.���@��EAt���n�G�<��祫���g߭��Y�+N�Q�'��mi ���i�85F\A?�qj}V_,��z���¤�l@�0�fw�I8g�xs�Hky=����eIe��m�귡�@�7��CD��ݢ	�_��������Lb��������qS*��kٶ�"��b4�b��*4��Ӧ�utږ��d��\�)dPI�fZ�kG���?~�N�����8��n�#I?L�m��9)*�\�u�4p�:��Ujh����}=�&����}L|��� ²K�G��ټ��h�Y�R��y	��߮Ү�s=�|��� ?P�I�0ɫ��O<�x��|�Z��G:��T�+�-�>i�Ѽc���D�����͒G덁�I�bW0�8�xY�_���-&��%S�[�ru�'�9��<<r��7����T�R���1�=�6�݈f�M��������#&�.f��ߎ�@�&��m-�%���~R���8���_���:��2Z�Cjn.�NO���邎����IN��tE;���k�)®�=��U�����G�RZ�ܪ�%�0��1�x�RP-�"�{\%�T� 
H�95�/�B4��fc%a;w�s���Y�� ����n�M�]�O.C%�?��ʔ��l]� ,�s�M?�E��?ׂ�-��*dC��IPF�
����9a�{޳G�����t���V�S>ږ(>�I��N�2� E�Tj���K�o���r�����#�mm軽����)<U�������iN|�es��z�yA����I%���ψ%��+��U4�0��q��(UtC"�Z�X[��C�g�`�"`��C�6'|շ뻱zP!`�N�3�`�Ā4�"!Sxx\#��Qr]S�ܭ߁O���e�3�/��>�0�zzq�� �S�׾n�c4�`�-���0�. 2�(��W�y�5���tU��RZ���N�Ee5Ya�KH�22d�{��t�L��Ⴢ`ɑ[W��h
�����;F?���F}���cŽ�qI�ѻ��1���Y�$�I/B`���1�n�@4Rr(�����,�K:�$��ad�����ɀ4[�����p��Yj�9_�4�Ol��L��j�b�ە5c!��%�Ǚ
���n>��OM`Vq��`��7�`�uw��U�@�}��c�:�r̼�l���/��y�ʉf-g1���3�����HY��ߟ!g������X�aԿ��$-F���o��j�ǈ�{$��H}�'<f��oĽ^��L����O�ijx���Ces�����Ǵ��7G)zKn{`��g4�p����� �f5�hR���Ԙ����OIj/�g�Ђ���snX7r^�)WCf��u��-���o�6��Co��s��O��5�5��(u�}��-�W� X�����6="����q+4._����+H⹈r�% ����׻��k�6�w�țv?�\ti>	�o�����z;��zX	25�ܝ�na�Ј�f?l���} ��+�-���i�Q@O�)�$D<KLE���T��Q�������`NM	ٕ��V|�{i�&7�cn<h���f8�L�8F�X�/��7�2,�3�9N�::o=9�iL��󓊥)���!�G0�����	�Չ`y��?� �>h`�� b��M�5B��>�S�Ox�_������ͶuG���Pz������7�?��?�,�������I^���	��Tnǉ�p@���kry������H/�pa�G�l��4����}�cxH��{)�u�z\�㒑��Rw�b3l�O�#�Y�w3�a��н��iA���#��%t4F���A�e����[ק�������R�{##������ɧ�P�PXd�����h-O6[��b�`����u�y��G[A���\����KIx��7s��A]^�_c���E~s���~;w�?�0
���}�u~�16�D����J�bC��ϛ�1����I�C#AO�t.������'�����1Fj*F.�h�*O��*c�Mvi�}����d���Fo�׻1T?��8F!�.󑧲��y��1���Ɨ�H0�?Yyi��k!jH<���5�\��ĵ^;��#�: ��Rn�Nc�Q�` I?�?�\Z�J�2ܼ��=�j���������%����N�{�FR���h̦���H��l�"�.Q�)һ��7��������yG���ή0u�4�"�S8���ΩS�J���y<����ʶ���%e�*u8D�&!J�9��LD٤9RR/���Fg��]�����ХE�v��>����
�1"���'�;&����jyN	���W��D`�l2�]��'_8��1/٦2er<��ȿ�%��E��U�����a�4�j���k_�%�w�;?�Nm��q���&�v�>�?Xħ�kv˦��D��%�ܚ��}�C�4�M]���;��5ш#�t6��j�.O��s�}&k�ob�+%��y�x��/]x`8^���M�!����?U�=��c�/:������ØUH� uڋ/����x6��H������W�>i��w:25�_x�^j����Lj���V��)(��´P�ǿO�v�ڦ��d����]���P��C�Jx��A����%�M���j�5�<�ʐIq	#Rsd��Y �2#�a�V#x�x@�����7 Z�s(D2)��9i��1��`�1U��`���	�o�TXD����HDxhbJbB<���פ�`7�Q~�g~���DǆЬ���C���'1$|@�T�4r�'^��E���
��ow�pq"e��2J O�z%����ܢ[�di�LK�p�eqp��)���y�2��{�Y��f)YV7�I���|S �0�T��V��y:;H�_~�d�lx��l����'����'в"�R|з�9����K_��4K���4:�mY��.}Ggg�js��Q�y��H���0}'�M*��q��p�+c_�L���s��A{������GJ~ZeB��k�����4��:6��w�����iy�Xz>��X��7���b�5��o�y�b�d�y��s������U���)�ǚ����J�o뗄��K�&�1^ ���?�\9}G�JsU�����@[��*P�(WR/Vx��s��AL�cW��sM:��ܧ/����}�pL`6l_��щ�pqa'&���~p���׀H��YI�bŕ�z���g�i�˽�����/|Y��Z\����1n,5dOrW�j�<{MZ�3�&^�!�!s�s�aPr\��yo(�w�#y(�[�/sЗp�����#B�C�ĭM�AJPh��H$W�̯�j(4�+4@�B,�2�Yf��k~�>����X0��ts��w%�&� �0�J��ĭ����y%$=�r��. Hre��X���ȑ&�+������ߵN<�F9��[e�J$�*�L�..U	�f^�N�����.�$.Ɔ�qq�nk���P٦���4���"K��f�03�,Ja��h��$#1�f,�5#t��� �_����I�����F�������퓯)O�^�ޮK@��@?�+��#����)�*#���Ir�|��O���f3��-�O�1[�����ʣ�q�^{��U�M<T����"6چ��A0�Sd�ӧt{��+K�a��S�����_\*9u|)�_�\s�{t� �^�K�\���q2�����ޙF���S�L�`�"�V ?0�-���G�aN�LS;sRh�L@������>����CK*���.��Sf�\�+(�}��
���m9�(#�-#@��-�iC��/�jȺ��뱵�j��)���O�0���'6ݲ)�TʴT!>�e�);���ސzh�H@%r��U}��I-"�A��$v�����L��.b��a~j���̕��Y�$@����9M�-����LH�Jh���m�D6��Kj o�������	z�7X2*)����t�Ҋ��[�8j6�n~?]��& f�:�0߄#+]�}��l+������Ig��tBJ2����ܪ~��J{�\��W�ܯ�녿���Ј?�,�<���ÇY_rs��؜�Ǘ37G۽H�X�?�ň��{�)���ƺ�%�k�C��b�:�)x�����WW�i�BN�)����!���%F <�����B&Q.4�~ƾ���JU�nS{�5N��͒P܉��u�nB�R'!t>��6@��a�6r#�f���C�G�����]�Б)�Ǚd�2���Sw?�>X>��p���u���Kt�Ol�gY�2�����݀�t��Y�R2y�$����l�lWW�3��S�@X��c���m
k�������UGv��I��':̢��Y79��F���t:`莞�iM��X�Y�9�֜���-4��O���<�qYW^D�+�3Ma)�?��pȻ=�V���POy�5����+e����l���Jޓ#b��vrC��մ�������z�l�v�6���|6�=��7=���eWa���t�ª �5�H�!������M̓������W
(�<��+�m���X��׊�0&�޷k�=F4BA ۳1� B�]�����Ɗ�U4+�L�D���VB�	����@�Әx�����RB�z1��޺����(�ۛXѦ#��V!�����B����\����
5���r��LS6F^�|� ��K�"K%�F%(���f�%�Gi~�|��P���Ŕ\K�TӁI�T}�k�H�WR-B����.��l��C���d��?/�d�h����(u�
m*vv��/�&$@7��E+���/"��3��r��|r�4b-5 �{�5Z&p��Xb��M}t`*:���.�.���YI3�h�ټH.*{n`f^UK�ծ,Ӿ!�B��bGxXf%��[`ß����9��yF�ϯ����ჄB6��$"�ȃR�]�[eP��J_��_y�8B�G���$���ĉ1K��#�+Q��z �-�`i��,����ΕoXl���������x���W�!C�99���y�����=�1�+VUQ�1��I����������b;�w�xM�B�i��)?�.*��{oզ��x�A8�E��AH8e�G�n�^[	�ȯ�ü�"|�fx\���t|Ƿi
�k�k��~C����{��5{�I*|��������͜v���Ж��y��ޑ��e���u<rCn5��=����5m=��_}mBrU��5��_syt�X�6���@yi��jl�igS.�ɑ���ʠL�dB��oh�=k�EW4lV���ʣf�9��U�B
d���,�� ��h���T�߼S�*q���D01�kn�z���,0�.��M
U1���$B:��G�q߯�*��o_O�	y���.����/%�ݕ;�}m�Q#��gO�D<�k0�O�t�Z��^Z��->�&&�(�1��)�!�/���l�d
�Rx(i�[�>cU~��>�/��h%�%	�C3�j���5�������q��|}i�i�Z�Ov�����%��] ��J��{�D�7��黤{&b��v�{�s�H��c�-q$������gtHw�g��=b�f��J�I��������A�;�MoZ�J�On\$���Dc�֬�W' �Ĉc���)˦N�[~�& !4��R�X��c��@z�X=}�:���7�b�m|FBv�����cr~&�W���?��=H��^����s��U�Y\���z�X����o`�	b��8/���J�*T��M֊A�ed
��FD@f����RH�e8{��=�1c�^*�nQ��&U�<�� !4g:Z�>D`y�*PC;�z��S&
G#� NI~�	����C	�oCT@%Qo�<ü;����!��	���*Ҋu�n"�O����d$@r�/!�S�����G>���?�l�	*+=]
��ç]���?r ��p�8\��T��~�y���C"v�����������r���R#�����%Z?ˊD	��pw��Wcg�1p/��e��o��n$KdkY�bޠ�k���ӟ],gV�5<������ɇ��u�O�/^�cl=��s����L�K�K}�q:�6֒ތCq���o%�I5iA��J��d��0Y6UgӰ����zA���-���`�|�� A>zY�{�F��)�ݖ�o��)��׷�Bq)k�{j
{N�{�;�nxd������( >űeR�lW`g��],��۴��1J:��S̎MܳP���.��%�..���^	C�9�D�{*�$:�7��1�O�м�{!�
VM�I��:����٘��2N�/2��ǀ���YAg!`C,#' �]�˗���6-Qȫ	8t�RR��eS�z;�J$���'4pw�(�V�r��A������um��MjbͿ����X�%'�(J�7&��l�{o}�#ePeg�9�S/hچe�j�eL��}aF��o*����ӯ��t]�sAhh@��˷�ɬcp�X�lƁ�ǜ����e���r��p�ƵX�R��6Ȍ�RW��{�1���(��Bh�]�G5�͌��z 7Ej�!�w�k}E����|�؏pzS�d�J�P�s���ӌ����������/���S�ݘ�XL+'�%ĩ���r�8�v���S���n�>_�k�\>-݄��^� ��{�v/jI�_�dQ���)��S����i��7����wO�W|���o�^��*^�	�4���B��>HW�4�>E�������O�*ĝ��E(�l�n��I��y��2��S��u�V=�$�J��Y�f��C葈jB!�Xݩ����ڃ����][՛�K��Pjs��'!VŐ �+7G�܌���'䔉M$fS��$"C��m�8ŏ[�'�q]`�[	�:s��{�u�sK{~փ�&r��n~S%�Qv�GZ��ɶ���^��k�A�`9f3��(9�f�SQk����F��^a�=�f͞*F9�Ȥ���z�H�7J��¨ �A����#G�s�J!���$g��bO|�t�|�VQ��p� ��������\2�@�o����Z瑫����%-V�rDb̸��t��8�e�7k�D�s&Ao�����	y���sF����q�U��>rU`�@�=g��s�؊]"��ӷL��&K"�3h��fF���dH�g�I�#V��\�q
��gN�>#z�G�w41u����m]��0Ν/��	gq2�	�_�V-v�<<�R�rM��!�������T�n4f�S���, �?ݣH��(�eo�T,Ф�G��|A�@,A�2Hc�$��rX�BUQ�&�������#�Zei�����Vѩ��\KP�Z�l{&Eq�f�Uƛ7��xVP���0��@����(��6q�1�;Z��tǚ˝��Q$Jl���L��z#׮�=��Z�4H��l_�:�r�����Wje�?{��C��5��Ҡ�	ihfU����
F/���A
5�h���Z��J�rS���E�6�~�|�f���Ũ��N~T�����w�Oo�9���@��~"����j�+Nzm�ׂ�)?p�T;-�'�2;)TM�k�عC�m���ZL��[m ��;�o�=�5%�X�<hR�<$�ck��]|`�!�e8��w�j�bYK���R�ԁ�=/��j�y4�&L6�3�P��W��#����]��M�<ޭ�g�n��)�Aq9p
��Ъ+�ϟ�A<�i�󨙛r�%o9z#�G�D^��k
�	�b��Raa���B.���+r��,yZs�!�3и��ސ�a/L��\��Nx h���캫�&��=e�s��M��Q�̓�׿��2�~~-p>&Sg!E�|��iE�)+[gw�K�HoaT�K��LNO����F�%���D�����N�2c�glt�:����I��K����ꊜ�Hau�ŅӍ�m�o�{f�,&�	��D���	�X��Ȓ�Iυj�vO�j�}��j8��:0Aྡ�Z�h���2���.�a����|��o\!�4>MR�G)���R��?�=ϥ�f�q��&/z=O�� pZ��W9/"F�r	�S���VBcC~��}]���WJ��yŵΛU�s�zЊ� �BGG�Z6yn\��&.��A?�qn|�7��� ��i?H���>�C�k"1�m�V�Y��~�����@���'���XL& i�g�
}W�Zb[9��?J�(���ۇ��������?���
bQ/� a�_�9Y���c
�n�����TF�6�&l7ѣ�P�+�F�?2 11�ρ鳿>>x>��:L\\��ئ�/�2�{c�K'S�!����q�o��VBz=N�'��.r��+l�"�k����?@�(���X=Ƚ�����a������{^�`X1GD�*�b0R���N�?� ���eR��Dk�s�� rj��������_��s�����h}ɡg��� �u+I�u>�h���A�1j�u7t)�_��mol~������r�o({�J>�W�`��}-�KaŤm��es�a	r�g�7�
_�X��ɫ�{r���:�x �5<��I�����6��/x�V��F�Kh\����Igu3�n�T�.��������.d�����m���-ݿ�hJzj d2��n��Ԁ�"�O��"�ɋp��gc]iy� �ܫ�A�?���E^O� *Qk�߈��&Q��kS���w��- )w�bl��0}?X 1�`��}��~D�P�"i	�l��0N`���m��P��7��o��k�')?��9�-��+�]w�}C"&K����\;& o�w�����Οc댇c���u'F���Vs@N0�A���^t� �9���؝&��|g���g �����.���;.l�or)ǘ�?�aUy�U��׻������	�\8�G�e�w�3�\bXL7(7�ݰ��_��%T��7���DBA�Y~O6��P�Arc"V��r�Xb� ����3p�$z��t��n�;��F̂�.i[���Yv���kK�u~��l���̖;p��w��#�n&�ۑ-����Xw���<��EI��{.����L:w	���d�݂-p�s�PX.�~�T#�gB��aC���F3�I������7�x���ѩk�� r�����|�Rg���ll�uJS<q�-G��m<,$��y�i���er�@%sTCc�(���;��8�'U�}1�9_��{px�X���r��Ȧf��MKRL*�.~�>�qu|��}��^��ӌr�"���i����O�C: ����N!�%"G�q��0EԆme��fB�(�y�r���dg�C��z��T�+Y�oia�+�=�<���/��8v>aA�IU�3C3�s��^⯹~˙w��~
�3�iB?�^���-�M��������+���������U���IF�O�.���?���6�3ቿۿw��.�qչa�i��$�70�?�,{[G��î�'�����ƍ�/�9��&1U<�N!�:{:q+�� ���;��|��F-w�8чZ�vߛ	V�؅�dd)�(��(j}}�w��.����+��BY���ٲ`�I�c]<�z�.f[^:��I��&�d�{�s�}��JqW�W�[D.W%~���I"&�ą�@ً��x�����{J2T;���Vy�h3!����մ��c�c3���v>%3#j�j� ��/RBR�%��r�R���]���R���o���on)\�,�Se�W-�u�vzD���?�C	�W�����ٔ
����ȼ����MT?j6�Y4���nP_e�;T�u�@�Q��sݯ��A�B^��9�?"�NW�*DЇO/���Y3aڛ{����j� �����0� 8�ptGX�Ij~�v/и>=�����h_*����=9h��Xa��0�aF'�d��숫�<a�uv]��f8���sv���%V��h��(�R[�x/�n��n�]��V::�=�ͧ`)���(�V������i���n�����m<frn�R��ˏ;��6~D�r����pk� IW�6d_�	%j^��������j��r�?SE?���Z��z��_ڿ:����=߫�%���=��p(��CU2��Lp0hT�BK�}��P���D^�Ӌ�ŕ�D��Q����m-�G$�=���w��bghv���I�������`��~0��ͷ�e�UEuU�;[��+�˚;���őZ��4���?7����?�E��8��`�s���b���qJ�9%A�K����u���S�X�&s�j�qW�k�R�T��<��4�8� �3�b�m�����f7螩�\��?�fJnC�+�S�fO�"#��Fw�_;}�~��A����)N���s�+ ��Iʵ��N��C�1!��e�H~j�����3IT���)�����0��I��2w�.8]ȝp|�=�kC��j#dp�\��������v��r �*$U��6ҁ�>M�����Wyt!��[���IWts?\����|��c��ik�p�)�F G��J�qz�'����o������ �Z(�y<�D#Y��΀���Wd��@����C����+�S������NlGϕ����1�G��A���v0ii��.�zW��,�lN�o^�T�n"�yQ?�����N�i�Dל�:z)<I�O�G��f{�3���K�������1���V8�z��&t��ᰓa0Y.��.�&�VYl3��y�(���ii{�rِ
E�{��\Z(�sɝ��
C]��g�:[����f����� ����*��>1�^A�K
I��ݻ�U�/$�H��$��1�ex5#�yO"�Qkٿ@j�鍂�|��p�}�Npkc������sQ�cKfv�gqZ�V�*�S9*t��m:9u�1�2/I��f2��!wE���$j�ﭾ��(��_{ת@Z�S�L���n ���mw�N*�u^ڒ'�$#�����aj��wV��'Fɟ#�t���O��^f�I�4�<��y6�_��}3<[����wrД�`M��]&$����,{��k{�Cv�ϳ�[�O�l�8�xMA2Âl�>��HQZ>��ӣ��]~��o�$���4Mi�8�웎dO����l���LXD�����q��\e4���$�˹��E�!�(h)�_f0��^/�.�t+B4O��2����Z�>o2��Q��ʯ�-�FC��lA�J(�� g���&�WS�L9aݪ�$g���̓�i���G7����g�2G����<��T;�x٧.i�_,'�����![צ3�q�\bUa���L.�+Ɔƪ�!�)���Q����]�oz:��jx���ۣ��9�������p����G'��-:+6~	6������(����`J�zf=u?�;��2� ��Q�}r�f ���W�MCzzӬ�a�n�v�Ü��t���Ӯ�T\�]t�q#o]���Ryĵ�&gǤ�]6�G�+��"37_���иleƌ~���4KIQ�����.�P�*��"�(_��4t���M��������+S'�S�Zs~>��XD�f����v�c��1���qF �x����B@��1�PI�Q�5��k2#ȴG:|��x�6��v�ԧ[�16�N7����GY���YYS�B�C֡u��=1UC��y٢/t��k^�?�7|G��_0]$�V��`.#��gu,�W����#SS)�������ڗ��C�8,?���Wx\a���YD�ݏ[e��3U~�g�M��7r}�K��6�-46VT�>��@�����[���̜�ݫ"����WbvV^����޲���	c�� D��o�
A��~��[�w��W���rSg�ߘ"�Des��|�A��h�q}��7�Y�eh\3��t��k~k���,iY��B��h&@�7�w�C�O��~>������~�5�l ��$P��SĪy*��� ��@��B�J++9F4���`X	����J����l����b
�f˲�8\�债f?"���>h��˹^"��IN-7�AQP��Ԣ5����XR==y�efR{'�j�/�AƕȄL�P��װu���b����룓A��r���"޲�{t�%�����!ٸ0(������}ߕ)WV���k�[%ӃN<9N[3Xt���/0>�/I��y!�!�e���;��!�G�0�h�)b '
%(ٖYf�HU�M��b�b'�]"�k��
>Q�	"#��P�[�z�ӂۖU�~Q�H������(=���ƸT�����������$o���㧟[*���X�6	���K�ۆ7��+Y����37l���lY��=�� ���(գ_y(�������o�}�{�V�����N�h�b7�/�ɣc/u�J	S5z���=���� ��Q�i&�J����w���D�3��(�r���E?IF�g�RY`�I���mjT��'���;��y����}�9���Q1�r*{�0W���+��5a �G8��A֜�4�]�[����p}�}J�@��c����$+���!�G$�P�t�eX���-��܂��Kp'�;����@����.Cp���]>��s�w�}��5?��g��j��Z�WO�5���b��&t���$,e�~�����ogxI���T��gJsG�� �f���̾�EG���I�Z���Z�T_2�ꖶ���4���0#�f�$�a~#��cQ?�����^����\9�c�aH�D=DJ�>��j�����vc�R��2DJ�G��sfb����:T��J����>j����)�^�����P^I��{�mx��j�QwH����ȉ]ͪ�(� ���C�v��Ǎ��]n�k��0[9f���Z��d��埽Z�|��#5�c�|�QTr�ӹw|0 �pZ+��^�ɃF�V|+a���[��q�v��;�����Y��bE��j%���f�}��+�js[0x�D|�~�s���Чk��_���1�|���1J�#B���nAR�ٞd<A#'��Ρ*�������@T��و^qK�L���J�r\�9tj@����ƿ��AC�A�!-������#d��\��¶?J_N�Ju��@dd����
6H~H������ư���ch�U�)��p/5[=C�~=���*&Q������`�/�_���d������f��!��Ø%�s�n�%w�3�[����X�,����Z�f�.Xu�ݺg��aL:���8"���P�?c����5�D��w�t��.�����5���5�k �y-����>���y���^��݋^��$�?�j�X9"�Ui#�]0~��0���e����B�HAz�ua%�x�j��bs�0孭ȿ��UF��7�����___s9��� �A%�uU�c���@������iZ�ry�wK��a!�G�d��[��A�yJ��[M�>��`WW����m0�e_-m��U����a�����ѝ�u߽���.��ɗ6�ju�y=\%\*;��c��ӟ���/A���\TzH��/�ޜs��w��B�/Y�9qN��+��Q2?��7���3�gd�RH57�G̠�~�m��쿯�
*�[�c�c�U�D�'���:��E��ȂQ)~�`܀=�J/�%9^��¿GLB���_����3'����bO导��zx��%��]�_㠺�Z�X����@�~Fbյ���ʃJY5�k<�oX�˃k�4�}b�
�����,�0@ԛ����EL9�������e_ƿ��8��(^J(Ю�_� ���q[-�[�?��}�I�[�p�\�����7���G��m�N�����x)c��uL��>��-^��J��e�쿌@�NyI2���ň�������||B���>*!V�n������sN2��^��\U���F0��BjK-Va]��n�	������&y9ܾ-�/�K�`rrϯ��@�RYȆ1.�~"��?�c;69g��PR��4%�?�B�bc���\���$
�O�K�Z[�l��ʌ[q3���s��@e�/f���j9���Z�C�XN2���9[KKK�"9�Hy5b�
 ,R� ��[_ŋV�����7$�]�_ux�������{@=�a�&O`x�#g�| Q���P��e@-�Uu�����nǣ���=w������2��`h�U+���g�B�
��D�)͞����)^zĩQ;��W	ߘ����)p�#��+��h2��y�a�h���9$p�K������%�تaX"����y#���i�0�W=1��ڥ�k�(1uJЈ�?Og����yZ�9=��a@d0Si��)J�#��_����(R��H���*� S�g�\s+d��
л9�:��Ka傿h�O��%D]���2!%�'��0�Yϔ0@����RM���&�s�\����ai�+[��:ٿl	���o��)��iF/ֹ~�ֽ�F�/�t`l��f)�!��]���pR�&Pw���*X�4���|9GF�_��@9�	iq�m�x��7��e����d��[��@�zҘ�5�W��}�l�7<y��H�^t�O���qm�b"�0K�Ť�u7Jip�U������%`̡�/M-J��x��\��LH�l=�Ey��:u@�A�k��xIs�Z�;�y{fwօ`�')���}�����ҕI��x�[b�
�2B�Xu�����Q�T��U�.��^�n�p��~�_��B�#�C�'3��r�q�$�� �Yz�n7a�{=3�7���,�Q�M��b�#ƅ#?������<0ZT�Q"��f��P��c,f��t�30��eD1q	@�R8]�'Q�"���8�gI�b������{��]
�i��7�ĔZ��>h�;���J>��^g���'''�B��5qqq�NNw�����a�f7����X���˚2���x��,('l��]���-�k��(�'��
�����-�I�aZ�C&�~����J�[��8�w�ω}���I�h��g��y�!�cV���QD"u&dD�(eu�r")�&|�v�?���ZkO?��?lzL��t,�L�k���Ҧ�*��ZNpX���������Y��35 qȪ&(8%��X���z����s�7"���=�L�h�j��Gv��z�*IOx���_&���_�����xY��|�r"���1���C�+`u����!�/�8AV2O%{ �)�J
_�ڰ�?�Z�QG9�k4_T�Hh�G�`��v.���c�� 8y2^��f��TPf��z$�-8ur���L���ͷ �lj z��{4���W7�����r^�
5�I��Cfj��Y�s�pj|d�����S^��b�!��7K��L�B�_������h�<�t��E���΃��zIGrME@|���Kc��U{/��~\J�&��7�;����$��N�.��̺eu�&cq�nBFZ�`�a^��ыc�U�/h)O-��a�ң�pR�}o�1bp���q�1�O#���:�k��q���{�����4U��*|i�� �xd|bj找����BMA�B�߱AT��<Ve\4���e�4��_�O�kF�E�P�3�?��,����iyE�5\�a<Pj���\���8��5�I������ϻ�i8�'�����,ׂ��t�E�������{+����s^���0�1�~k��V���D�i.�s�w�b#
p��7�g��|T�h⥮me ԁѲ�<�/�T���m���n�^L�������>eb�C���K�ʲ����l01P#� ���"�U��O����*�hT�'�h�̗�Xa�@�GN���T`�w	�*�~}�"7:1"J �͆:����	gK!��vy0���=���+����;�[/
Z�S�^-�1m�� % |�bͰvl!7Z`����(��-f�0�:a�����*�}V��;}��>��E^�8v.#'*X���gl���iҧ�f���ŭp�!"�t�L�[��6�Vn�gT����?7��R�V
��îqv5_���Q�>��ZJ<�Wb��N0�GG���څ���1Im�~d�՚k!�g|i�7L9��h!�*[�c�l�;ۻif"��^C���jA��^�Dt3m�>_�,2���@3n���$�����\��DD�����E���=���X�B`:�$ �^�˶�]��8���/#W-�Z˄�&˄��`��F��uי��U�+���|�J���]1*ͧCG+m�?�Xj�:��ǵ��5�`;�v䘱�qXs�i�
�6��������������U��CrJ+�h�#��Ҏ��3~ˋ�c"�lf�͜P��dy�$m
^��`#I,X0�Wn����\w��F4V2��݅��_�}�Xi�`(y�i$�[i �{r�+wl�߭��3yt���p���B���*����7��.zڤ���w�d��ݏ%dJ��ŵy�E�l��̷(}~�7�f����{f�����-��HNϾ	x���K6)2���M��4��yإ�3��7U8���W$
(7Z�ݚ���:���+�ח˿���כx���{^XJ����O�f���~�AT-�hLʷ&J�t���?3�/�&�����D4��au�!l��4�GC>#��s��v��G�<�r4��t�o�.�"�K��|��ټ��������V.��M<.������D�E�A}��vb%~;���i���M�7����Lo����ճ\��i�8�]����呢�S�=�_�ti��%�'�Ag7e�|�{�4���~TZ�L�k�Y���C��g7liI�cR��PV`�_��!��N��7���ހk�������j�%1q�Č�~jO&�~�+|D��t�#��O|w�3.z��fFѯ���?Xft�e<I�롬���&�uʎD�� -cɂ,(�`�3����J�;j�Y�IS��*k��ȕh���F�u��O4�iXn�O�c���R���F����r{y�a[�~@�������х��UѶ@$K�Tۓ��,�ܚ)X��ѱIuU-{���_q�K�[hߪ+����'=�b���d�S��G2Ь��F�����:S��^�F4nz�y"��&D��fg�`�u%��=��3tρ-[��~��:�G��D-0;4[jB>���[�h���jTi6��)�K)���g��q;,�Y�2od>_������n��,Sp���N9���¡�90N{zEz�5H I�V���Np,�P3׫?�?ldB��
6�vs����?H�U��?��dS��1@D����}D��X��Xx�x��x7Y�R��/˄�3�+U�"�R~bd���7�@�$�����i�x.j����_٬|�i�"�Ϊ�`lA<� A�<�i?J��±\M?k���)k��2�;0^�H�hI>�9=4���u��L�,��ʶ'�6�~��ŧ����6�4{�7�]�_���D%׏ʑJ�[
er�*
����Lx�z�����n�t�KD�zr��ݙ��f?Q>�
c%�9w=#P�"$���������P�Jm�}�Z�k���L�W3lE�sMarԐ"�?�` 5`v�kVq��3)<?'�!KR��/ݱ�˝?R�çݫ��~����k�ٶ:D��S="H��쁤K��ḭ�]:��/���O?Mn���W���)L��FL�&��Fl�29,3©����,��uп��M��*��+�~=�Y�+�F��۝���v��~�`�̺�,���P	ʿ�I�l"�pA��6]9*���6���);�٬쉵%]��w�n��{x���=vw+�o���OҶq��a7S%����Ѩ�	�.V�z��D7����6��-Lz��L8 �]i����r��&����z��<�R��J����?E�����@�)�ԝ%�N��қ��ʴtZa��,�?ucZ��`���^};�Q�^����~�~h�N�����A<�c|���<?f�4�Zi�(�<�V����z-�N.����*��閗(7�(Ugܟ��X�U�<����t�[(���H����4$j�q��-�~1�m��W��C�*٠p���&�+�LKέ����ߊ޽�
�`}�n+��o.����:b�60�4M'��yN]�F�҄��7!PJ�'!<���(uP���&B���Q�A	5�c���ft��a���`r�I��x��^��V;�_�+�ƴ�zH�/˫��î��ם���D\4f�1Vfe�=�'��v��Ի׸��LtC� �և���ʟy��(����Z�%��>��'+�LԸ��
G�D�r.{��_ߊ����A�����Q�*_�G886�6oTȌ����m��f��Gz��Em��欇�3����;��Q���6����"���p=��o�b0�ig����O7M�c�^��$i�;A���Ng{�ɑDJ*��_��P��k� ���b!z���莨/�q�M�N��p��i,Ƹ�\�Z��_�c�j�q�	�'L�^w�����Ɍ�����e��j�Dc��nS~�A��{d��Gt��@��"����J!�TZ^�Ug_z榔���n�՜�3���ߜ�ᯭ:	�5b~-�zrn�����5�{1���ǯ5t����W$���t�:Gѷ���F����e���a���k�<�	ޢB������?��L�m�}����U$��E���Y'R=���n2b�=�垼h�n������Z��G��Zb�Y{�h�Ӳ���j��� �2���0�Õǰc�C�<���"��1���~��-��N��J|�2!�Ä�D�(�QRRpC��� He.e]�mU�;x���s�(�L�[�3���Hԃ? E�͙�x`�K���k�c���Yr���q6gAQ�� �4o�qt��A~�Pt3��X��9�"U%��!~$&#���/���,��ّ���'+�/�����=6�ʽK�:���n����j�����b���J\�L��d����m�-��Fw���� ��j}[E��+��Y8u�/Ҳ��kz��i�X�p7v�Rц'(E<�~l�L�fy� <j��c��	�nh7͜�?��܊�{2�sf$ޜCͱx�����p.�\`uށ�Gb3�}����l��8H�s� ����R��JS�Ɠn������Y vd^���q�r@7��i06����_�Á'�6�����}m0�%��Y���6ID��3{QU����ޢkU{����F��ĵ��n=j��R��â�~"}1�d��n`�#�_��h)�ȅ
��lC	H�e~�v�3�q���7�vf��l���Z!��}Ҹa���D�W#Gq;'Vn���bsءf� j�ĳ}�6I^���ʃ��`N���8�q�� ���+P��s�W�jDxZ���Te4p�m����4�r<�Z��<�ʾl��(N�o�l�(�v�#h�d�UI�$)����ȯ)=���"aQ��"G��,xBNM.������`���i���?J"f���G�4a>e�;o'�[-ߒ�����鷙\f!#y���F��)�a���<�:B)���\��H0���g��gW<3����5�R��qH�} �z8���E7������.UA#'�<��Ò4���=/Oм��o1��Ԁ%g��̪�ᄸD�gd���5=������f�]�G^�-����,����V��nV�O���wz�nc��l�L�	�hk?녢z��׹��&��D\�<2���r�o[+.��D��y~�C?xG��I�p����l. ;�UG���;NU\��>�<���sC�Ĭ���Wm��Ɩ���^��=ɶP�-o�H^�S��ּ�������
����D�5�Z$��'�������%�cTQD�O�{u^ ����q�P�P6*}�d	��l ���7ѻ�c�
$��q���˂�����h1�']�
't�u�������-��uz��\H���]�����qATDC�X�#�V]���Ӵ��`��21 ���gC�MA<��]��ռ�5���%�����$jY�!
���	����FZ�P��0MB_���m��@^n���i��ŧ3s��V��Z ./E�M��HC3~3����;��r7� �V��%�^��Q�.�����K� cL�R�����@-a��D��'���sP2v��oG��.�~aΩ�"��D�Q�"�A8�<d�hl�xu�|�,�)y�Ƒa�;	4�M\�+�*V�A�%0�e_�_0�1P�5s��8��<�����Rl�Ɖ��4TǇ�ʞ�|��-Yv���6)���0�Ǧ��`-
��������U�3�ʱ�{`�	��&;=z������ϱ��9�"RD�nJ���u:�38�_�jT{�Wɠ����ZF�uI�s�`��'��d�aP 4��rKK�ǟ�یR�O� �>XyV��3�up���1P��I`��M��1�eB>*�-��_�({�ˮ�����z�ݼG7��z���:1�@�P�[�8�I�w�-<h�8�j��;p��)���¯X8�+��et�6�����Ȁs^�_�*�%R�mM�J��B��ML�v���<�x���*�4�mbs6}�O���uU�����б�橼@Kmh/[^vec18��S.�Q�7-��Ҵt��yn�\��D�� ��J{�Vq�H���:lHS��`��Ƥ�(Q�0Y�	�UIH�9C��}�#ۜ���Ӵ �{(����G���TM�33z�*Z�*Zx�櫊��%�vq�s���bߵ�z`���)��'���_�,��C��x�0�����H�:ar�%������׼@\����O>B�d�Tu�,�CJ�vxn�-�^O���*X�ob�2�����~W�����o�Qj��.W�M��Ϋ�##��9��ȀW2t-���ȿ����8��"d��$V��Ћ;��3�Jf|d���RΦ`eq@7�
�r2�{�M����� �J��4�.��H�n�@LP� ~Q���\���j>�G���jœ��8L��H3Z��T�W�h�9�8�b��e�rcdw�Z�KR_>7�A5�&�.n%%`�
m�mfS�+�M�B)K��E�T���wtw|�E��Æ��&�J})*�Wh83�Jtm�4dA����2����oP���:�ˣz�7f��:nMȰҼ&Î����ۺ(H�S����ΞY�=Ho�\�_R�L�q6���­��4, ٥rƴby:�3���>؞k�p���5�������`"R��a*Տ�ϭ�A��|FC�|���2���鍞aw��Z��Rya3��$�jARRږ��o��!g�⓰���w<��P/C��
�ՠ��'�^h�٫�'�pV6���=�[?ҵ�Z���G�CC�	0�6�jbj̈٨�
�3"�~ ��u[�s�)#˰�L�2Ϸ_�,N�!w�.wK�$)]����؅�?ë1{1Mw�;4l��t�^J��߂��[ ��~��涝1��Ϻ_�_#g�tx��+���^�}�?9�X�*[�<�~���:�A���K�Ï����T�!	�[\u����1_� G#zN��=�
l�?� R����:w��լ�L���,
���W������B����%-�k�m�j+$��v\<��HA�R	��}(��6�V�-	Js��@��;�j?��)��S_d�Q܈I�x�]�[�şV��/c`?�3��V���XQ�?j�P\r�Ų3�S�[��< ��­�[����XE�ֶ��F��R�,����UK球�gĎ]�����*A(.�k��T��.4������>�'
��r�����&����·"H�������o�j�8�`�!�����P�V��3��4�!echkr��:�QD���(�h ��s���C$�V�~MH����S�հS����ae[�ju!�JL�)O,۽��t������y+��({'Q�d$�=��سP������a+�O�>C�wz�&\�����^������l���	�mk�l���B�^�%Ӂ�>�(�-���#0��(�z�/(����J5�G��ܟ���Mm��X�z}}}����dT,�_MYW�!d�ޑ��WU�%��3q�1!"�>�xN�]�]*�Qv�[���$���Fw�b��e���/x�ӗ}��Dő"���酣t�}��c��-?��������@���g#�l0 F�S{�����w3 :k��i�DŇ�b�++ñR.���o.t|v8縒�^���1L�߆!�yxb�GL�	"�є4T1�Z������	�+�[���D���JN{q��_�4ΒF
�_�7;�����Tzu�m�~W������v@v� ���W/rܤ��a-�)^)�� �RL<�	\�J�\|r_G�O�X�bW@��2+�|�?=�x��¶?N������~�Q�cV"!s�>���N�M��u^p�뷞곕,aQ��>�7��Uq�\��[J�!&�(@���`^�/Á�����u�,�S,� -rh#�0����m�S�m�fM��׌3g�J���`#K3������#�^0�`���<��j�A4s���=��ͷ�>��/�[#?�#��D$!BL��Ġ�I&hf�Or�ԩ�$nm_n4��k�tc)&�['��ğ�C`�"'�Z0�{)�N��4�v����M	��h6�lX�|��U��� �q�GI��$�+�[��%ڪaX��̦z�t�/T?	!��a,A�����^�b�_�W�#�HB��f�7)^@������.n%@����P��,pV?3S�F�Q��9��8h�9q��h�?쒴�R�rDvTO/��Z##�'Yg�!k����8?��h>y[�5�Q�����_V� '������Ô�}+� FYta��v呸�X�)�z2��u#Iev�jc�X\v�B�G��`|;z^�0_O�J#
FbH�1ym�������
3j1���]�Z
_;���F�Mc�q�쉶T��A�����q�,��}����c��~��n��#��t{�E,�8�t;�1�����̯��A�<��X�> 
W�!�������vҢ�D�%*�����}��y�8���9���>v�~2d�Xd��h��Msg�.���e�H��=� ���D�h؍<�S�uѧ��8;�;�G�q$�^��X���B5f}�r��C��T�"�z��æQ�CD�|P���"| nQ	��h,�#/e�}��4N�/[��<iK�$%��m�@�����q�xD���?jd��[��`AB�uz�B�F����s��P�,r8+K�߰��2$��;C\TQ�2C��|�&#� ��~�Td�Pw7M�����c����VM�e�br�k3"�i��3��$�đ��jT���⺕O��p�J��.���e���S�w�`'�!��.�DKԲ.� *ӱ�4��f�#/P	�%�&]�l����:���N���0�ooT�����ǒ@,q�ɔfn%���s�>�'���en�ܯX��1J�<�ֺ'
?)NqR�$�Kz��O�ܬ�|�]�+�#\�
q�l"?����\��&���mj��T<'�?�5,_͕����D�<O�0�5�lW��F�	�P�H06�_W������;q���V��K!�����ͩQ�͐|Y��	F�WpI
n�*�g|)?��<��$�!�P�T��
w�.��2ܗ��ZB��\@s���#��Qc��7���d�Ms�f�����f��k���k�={�q�,H*ר����s���^���dKN�+���ǊBC�#W�P-����a�BptȼƫD��כ�ji�<%Nɨ��Y�i��pL%�D�{ƕ��`g�($)w"׼�)MD%~�������ne�A��6&�D>�t��7g��@��ue9"Zv���p��7"���#�� an��ka0�c�$� ��C-D�~(C���A�g�*��b)KR�Ӛ��~���G ���!9�&U7Q~_�ǻה�4�
~Ge*��O�hS�6�H�+q�QF9�XP� ��'2�\Sld����w l�z���X�w�o��a��Ցq�2i�WR<��4�ݲ���dT��j93;�Q�����,�&j�#ޒr����Q��|J�V��a����09^�=܁r���������ݡ�{پ1��0�o8ԽRo�R�S�@B�#E�%�ʸ�!��/JqЀ���-��*���2�U�`�$��̷�)Tu�b��=D��ʚ�m�/��-_���	�E�|�0�Da����VzĻտ��TM�2�Tа���KA���fZ��Հ�Yg��̉��� :e=s�T����\�,�̂��D0o:�S[�k�Ff�v��1K���I��⍠]��e0h��d� 
D�R�v�|u6�e�����l�?�3�`AA��3\o��5��;��Hwoh�Ĳ�-G^=�m��'Jj�
l�����h�����e��h-q(#i�N L����=y���&w�'�C��w�߸˱�ʱ�܆�=�|2hƧ�*M�w�Ҷ�1w�O���D��/ 3^�x���s����L��4d�Mt�#L=�l�(����x$�p���M�Ƶ>EȎP7��^�9�A�-e+�U���������>E"am�T��u_���t�yh�u�b���
b��U��	�����I���8�x�,+^� �����Т�� g& �
��i�s�j<����?��� @�Y���_"����hⲈY�d ���r���(���8 ���y��eʸVl�MhK�%��k�>�D.d]��c��E=�����=xw��IߧO�,�ysk�͋�
�2W�5�4ʮH��;�1�Oއ�� ҏ%Rq�W�,�Lo�9�gkǾ�,��W�I��Ci�\�ڏ�q룙X�bi��D��[K��r-2R������$�F��%�I�F}�i~(f/�2�2W�:���e8��1r:�����2��M�R�1�T�ź!����W��=�S��6(�2{4k��4�{������ }X�]��;����N���A=�����_^��Ii����N�߈<�l]L�]���C�c�%W�;IK�i��`�~x�"&�=��=�7���G�y?R�)y�~Ijjr��do�%W1�(E�r��,M��p^I�pN�wCy�-�:�7�k.V����ܐ��O��%�O������]���/!c\�/�5l5�x8)U�eyF-�ᓏ��/�����e5�����Ы�a	��9����.f � I�PsV�>�8E��$STW b� �T� 2T?]'/�%<ɤ���A�?z���\��m)����Hx*�n�)��#��[q��hS#C�̳D����� ��|�'d�?��[��h4�>��uK`�S(;����h���s'�#��bR�0��)�A���hCs��͹Dgm�zv��%�d�u��u�΂꯫6�g~�}?v�k���Rd]�o�_F^ck�C�o�Rn�Hy�U�Y��{Q|[2��Ν�	m���(��sm�?\���P�|S����:|�Q���Q���OW8�|�e�8f�=�H�vFh�����!Z�����ف��͒]��nQJۡIǐ��u0��#�E�w��s��"�R���v:�����=��я����Mt�w�Ƹ�ݺ���Z���<����Ԋ8�څ�t��:̈́`���u��Lgti)g�"�P�܁���A�(�����?5��wޗ/Mt;�SZR7T��ؼFQ!��Ii�Ӽ+L�Q��������%�Kk*8O�uQyඡ�� ߗ[�W�"��R@�m��g��SAm��FL�fNSb���T���F�	����^3ύ[�Kt����Qq���;�nl�28^'�U_LKęku�\:�h�S�a3r��R�mM��<�ho;���� 6�9sc��� �_����=���8x�L��~Ґ���>�¾��T�����VESc����5ژT�l>Ļ�=���E0ds�|�G�W�T?�=o��FWkG�����|^�d�D�_�4�5�M뚋�מ
��j�z*���:A�{�%of�/��qT� 2`A��sJQ+��Wɇ�Nږ��V{�!d��*%|Vv�M̙~*��*���[A�0��qF�h��_�LЧ�����IF�I��]���Á&�2tы�@eg���ʬ�_�s>m|�oH�M��o�\��a�8E�k3�g����~�kO�� ��R,kJe���hh�/Q]���뚯��	�l�zu/h�g�-ڴ�1+X��u�W�\�՗,�\ҷ���ݑ��e9M]gT/��xJ��;H�E5�r��z�Q��!�'oq-�B��]�l��9&]�NK����[���)t��s"��.�no=�zd+Zp�|�5r���q��=ט��$�m��ǩ�"����}�[J���9�`�.����ƲY���{?��n�g7��=���6���5�/_x̔z��ܤ�+=�4ί->;��f��O�-�&'���l3:ӹ�O��"���d�n��t�a7�O�z#�vH�|��D�FG��/�;��Y��F��:V[r�(���QW��� �I�����h�Q?�q��e��Ƃ~bIX��w��������ãE��7ˊ<�C�ǆR�q�#��jbmނ3����΋�|n��c!�VK(�&���J�lD�I?֚ԛe���q�=[�0#ىɖ����
�,S�1Q����tT��/jV�������$;X��g�{-�޷�e�t��y�C�~��Ղ�A.Y����<>v�ڠ���@r��+�2S��� Q׌��<4�#�M<�6���)�NȘ�$\`n�Q'ے�κ���ָ*ㅩ�K�%
�q??���T��(bo��o�� V7s0��:N�0��j�CGR�N��o� �<up�BQu%���+V1p�/٩�QUn:�y��
�?i8���!(�-�/TI߉��j,��$�� �t���l� i�n�}F*|`�����Ϥ�d�������|�Q��s{���HC1���c٨��C���x���Ǵ}��vWL\�i�Uj�������6��^�����J=�NϘh�P�N�䦦�+��zd���Ƒ�|��B>��۴��o�� �>�B�%�NSڑe���q(�e�8�}���pK rH�I!���	�727\�<;�;��ذJ!ij��p�je���=`�F��zZԌ��;��XQ)z��x�F�z�B�[De�;3g=�|k�#�.���n��}��߇k<�7+ M�My'Ԝf�
?_�`զ��� (Q�O~�=O\e7Q`���M�j*�K?�{k��%�s��m��WV�x������<+��Xp��6�2*=�y�M�q|I+�p�, ���*goQ-�>?���F=��� ��<���|�d6
VM��*�N�K�pĶ7�ؘ_��6����M?��{��x��;�yd�/^�4�	��Vt��Vo��\��	��d�lb�L�] ��Daa���;�n|V�L;zZc(��|�0BxJ7`�A=W�Jg��/]~�VDXty�5�?�}Q�@�Y}������H���R�]�T��Q]��ўTݸ<���qEԿ��謦�kgDre�3}~Ɩ\�-��t�P�%�5�b8��M*%�^� +����a}����=�-��c[v��r�d��5r���W�5���Qo%���\G'�M{>�*5��=v�Xs6wCc�3��bwВͮ�'�_
ѳ:	�����|@y����ᇹ�K�T�)��	��׵0"����ggW��F�#�_���+x����(��(@�V���2�_-���M��q�q��.�0�\��vKvv9q��_���9�&�B�SOV,1����VT'�{OOA�zQ5l�������)���R5G/4^�sOǺ��D8ajh;��?\)�v%�j�o+�/$���H���7L�֓���Y�7������"�K���7��1_uI�C��H�I���ue�z�	�����N��\%ݝ��s����L�z�jf������.z��Uw���Eo7o4�0�����H3z!H�S��qt�G������fJ3<�loE������.v߷[7bqj�Ie�a�e�r6t�A�3ܧ2�5�B�B>\�+\xk�Or��Jv�d��DP͗��?�O̼�Ѓ��px����ct@�A���c�\Z�����y�NI�vN�4�]��:�a9*�=��~���	�8�Ɯ��.��Z\t�@��$�9�����G��tn�s���}c��qZ���6�:|���
��� �*�
�n���H��$Ӛ(z�y|#�0�)�W�+7Mg8�)�K���EĀ���8|�)İb��CsR�� L�-���!�1ծe��[ /h��i��4�!�+MFO�BUr':�YiWc}j���"ޡ���q��w\�� K݋�Oׇ���̏��qu����cW�mn%��Pln��&: �Q��m��鰹w����G{oU��m;�1���y)0v0y'�h&��nufr8,���&h�bu�>�
����I"�{ۑ����r��)û�����ѻow�VG�ߺQ���kL�|��c8�Z����oɝ��g�Hch{����'>�Fy����F* ��N���oUW�l j��p����Q�]A>�]'��	e�������fE���Br��	+;����񤒤�*�F�����_��B�"G�|:��Z{�� =!sb�o���9�F�Н}@��k�換1B�Pn)�ċ�x$8�M�pﺓ���*�����D??��q�9z>w[��=����ֺ�R����
r�,l=�eF��1����λ�����џ���~�*��~�)<��U��Xu-����ͥx-7�s���Y���qT����Kw7Y��՘�ۼ}xR�#��b�~a!����:jp�2���b��� $��x*
~M<5,�@�ވ%�<�W�9��(�H�Y�4[�7�u�{����1#�e�UMG�{3���������H�Ϋ4n	������B�oso�1Q�p�Gag�]/��� "5e�7�Q�,G��]�k�
W�ңZB�/��J��Y�3�L�|k�g�>Jdಮ�P�^�U��.D�Җ�c����/|����,x�%��E|�_F�t�-�6 �=�7(T�A�����w�B���.N	bC�eK�Q�^Yv�ƶm�wl[kŶm;�������ض�1N���W�f>�T�WcV�5fP2bɜ^(~���	#m.�u��d�[�(c��Q�6�kz����V$q��[�oܒ���`�G��`=�����S�g���y�� ;]¸E�J�3]�m�s�]�ܻsS����C�����هb�kB��|x�DQP����k�U��ۘ�!3�f�� ���-v@]<���xK���c/`���w|9W��+,r�^�f���QAfY���8/Ȱ^�`�]��ksܘN��� K��e�_�5ǚ|?}t��/\E���b�P���/Y;v�$�Ђ�WZ���u'���� �1�k=�M�{ünx�OASE+v���iC�$C�[��NU��Уv��lB���0����=f�1�:��?l����M0���Y�����b�yy?չ!Q�G���!�b�	
x���u�>�|���,L8��.Y`�hR�"��Gr�A�Y֢��<M�٧�c�=�����oD�+���$dۓ��{G�*	B��!�~���v�e��ά$���&�8��Z��4X� f��I멄S���>��K�xm�����?*ȥ�����cC,N����Yc��
[��e�0p�o�c@�>��"�<A�fl^X�鷟�{��ּ,>P9�����u�<���E�T�_��D�����0��!�^�K҃����'n�T:b�+hQ�03�Q�h�12p�`��B?q�%h)�t�5�2b�b��p���|D��K<���H����" �~�6rq��ۯ�u��j�,)_��d�/N����V;��=�<uPG.|�t�q�wx���tT�^F��C4/Mi����3�l�ΰO(��|m��l1��'oj�]��z�A:|�p񉝈X�GP��Gc�I�8�s�ѷ�f�5�G���.H�28�#�û.�2�5�vʼ!<������D}O6�j'��0��?ϥ��,W�?
|���A���V@��er��$�D�5n}�?s��EW=�7�G�W�Y��ܙp���$����1����T+
�|!�_6ʡ��*�T�4���;o\��hC�#P=�p3�85�C�0�5K�u��}��|�c�.��G�I��Yα��Mv����RHGT�	��fSO6�c�REh�pF�Z4l��[�uQ};R})r����	n�j$_Њ|��!�Z�� Ć����0�h�սzG��A+��m-�RWq?D4�$�6�ڄ�1�r��JPү���������������,��z�������0���B\�v`�7�^S�@��u�����,X��9��%�d�qKcٽyh�+c�U�a+���-�҈�����9`�3&͐�����(�M��PC6�x���y�
�!I5��E�	�0�SAN?K�<�&�����Ѱ�͉��.�@��h�z�]�o�>��������?#8��n������y"aU��� 'L�ǟ��sq{4�-FP��m��G��WT3s{��0z�=�L���G�d�EB�S_�
�Vɘv�5��ߑ���h�x������\ T�G
J����
b>�B���h�֠b�b>6��z��h���ݭ�Grr���Y�֘y���]-���z�]nh�A�Q� `L1^��t�6K��]��}%�Z(c�qg-�=k>1�$�5�؆D�M[7&�
^o���͏���NuM����a��m�L�4�q+������܌��+	�C�H�\8DU�����VmwN��*2���R��м|�������Q��J��=t(���iD�L�i�f�c
�Hy�buh���wr\�lm�a؋=кI�BZ���2���
�°��/t��3={X��t��?��������Ifr�����[�MR�'J�zr��mLv��;�ÐX�q�Ex�/�뷍�'�]������V{�5*��]��j`k��$�{�ے�����=��O���B�MC���-�O��|#�y8l�	0���	� �������G��r3E|��L���\waK�Xg�����/���%Tķ��A>z��w��z����JLZ`���MN�@���e��Y��b#Dp�Z�l�,
W����,���`���Ӭ֊����sw�M�{�KOzW-x��z�~�TP�ݱ=��/�ƚu'���jr� �Ӄ�r7ڼgr�=�ǽ�~3�xGx����L�=��B�?�Z��r}k�O�\r1<����R�g��Zź�dH����3�0&oR�(
�xD(�wֿ	�%b}�g*�Ʉ��HGl,nǠoÎh[w���@:G�-k�h;ɀ���4<�>le�FXfj6U����>���*k/�VJ}�^|J��ag)�j�&t�f=[�ﬔ1t*��h�����6���<�[	�l��d�:�ɾ	sfX���u�К)���W$�YL��~f�"��Kz�{ٓ�W��0��U��b�������$�K�aі8�'Y�>�$�31�&rc{�ܷa,h�ر7)Y�
� ���^N��8Թ��!C��\��{���J9�VmD:�'�����N5b;� D�_�	�l叔�%A��tn&@#�˙����p�?�?�����H�������YJA?�BGyb�ڜ	<:�nc)6'�ޱ	�s+rh���j�B��Ƌ�]�<���$�-� 6/�張����i�;������ɥ1a@�%�lH{�.��׎`
�s�sQ��ld:7��M��6��1�akΙ�bO�	���G��y���/�S�bk���3��;�XRd�xU\`� �:�e��X��-�}�p�]X�Wo��ť��z����q��y����y�M4��AS���BX��O��x�*?�q-��*�0�[T>�)�����9�~�oŐ���/K��Mߞ�;?�v���������R7�����<,�}y���)��꥔�z�l��V�3�j�k�#l"�&��\�A�FBljvz�n��>"˖ dl�����%qXv���n;ٍ��D��j��#��/���
W��2����:��/_��W�_��T����Md ��z�%̟ M,�2*�ph��EJ�|�1�q� �꾓Ҝ������� ��P�ۛ��]9i[#����}��{tN��v���5����nbzn��F�R�e�~G���uCTN�H�Hy����ؚq��hl|M�c��,u;UT8s΁��f8O�b��e��}����JY[�����!fhF(��1y�����&�"n�i�O�у�#��	�o��Z"��Ay�4>dG����%�Rc���`�c'��B�B�{���ؾ}�}��[c�7|��$\H�iШ��-t$y�w���M��r�Jc��oM��b��Y�g�̞��^$��Pj�2��d��9�a�F���s�V*0gGx�vE0�8o������./�F��t�L���hq@�sw�}aͪ�����T{"�'�v��v7BkW�08D
�����f��e���@Ґ(	ź�##���	� ��Vau��"��b�V�(O�����`�:0��	���Q�g�y����Nt�]Xd q����d�$�8H>%���y�@X7�I�Rr%Ҩ���L{%�o�c��#j��O�%^szp�2�~���Y2�E���'<q�&����\$�#g��p@�d>bU�"�ƽ�3��x�j���ˎ��g�s�;�z��V���^�ށ��dd�>As|�z?���*v��}�6c��IHf�K�G
���+�?�ɘW*p��&''D�ٗ�ge���1�������}�S�)"R����w���P�⑜�>�`����;���m�=����z��N�1��<�z���_�&	C��RF�!J�U�1a�A�A�7N��:�I� !*R������۾W�'��
�	��݈�7��m�]���l�XD��`�b�O��=<f�*�pm�@���RR�y�^�z%o�޿��*�	X��N���}��}����({��8م��9Q��b��u��ӺT^g�6( fy�9�+L�5��/rb�|�~.?h	"��,�v�
�?t�Q�6)ȉ� n���nv�l Jd��V���ف!+E���&΁�a!|����EwBv�e�wP?��y�5;}�žlT�8|'	D.5���V�2���h����K������%̉�@��p�T�D6��
Xv�(��߶�0A R�B�3B �>�s���eSW�Hy�B׎g�#Dz}qJ���J(Y0P���f��i�AdY�.�Y�\��P����Ǻ:h|ۊ����f��
��/�&k�e�\<7�-������ƻ���
����[�5��x�{U! �O�?�j�!�b�mo\(��"������)�h��k����2;���:���YnFkc�*HM�Kw<�8�k��6���^�:�u򸈦�x�ހu��#���P��M�AA�6�6�)lHf��������_����h!x�`_�q��~���Ž�.���ά�]��1zԏ��Tv{�&j�"H��{a�Ks�W8wr�ND�s����5�7a��J�����ț0����3t;6���D�>5��I׃��h��S�'s-�/�*T�������~<BA���C�����?�5��ж��uO�lPN��5t9��B�;�&�͘��N)�Ԍ�R7�t�|eh~��:���]�p���g[K�T����W��O�W������}��yI����s|���o�����e5���ԉo�$&4������������F��B��sD���|nɓ��CF�*�
�S
7�E\�K��K�@p�Nu���UuN�W��N�������#�Cʁ=K��B�����|�Ar���~�;N�YU�:��t�?�qC���!���k0c�Hq��g�]���GKp������<fk��skvi�`:��j�jZ= #���3M�T�H�$ӎ�Mϐ�F�ܴ����.*u�c�� �ث,s����N���q�M<h3�`U}��ဓ�'�;c�Y<	y��H����Y6�f�X"�[X�+���ԐQ8��Zf�̸k���d�7�r(#�����D���GQ�� ��u���|}f����wi�4��ܿ�Y�p0ECcA��o������ɫ<t�by1�y���Y�J�"��(~/�z�]p��'�i4%m�w27���a=y�H�x��/�e�m���kfŜ��1����oa��qW�ku�w�ŀօ���ٰ�X�ޑi/��/2+��z��AD�;?�x�ij����ɡF$���Y�v\��{?��/̓��X�cn�;ﻦ�_`���#Rr�Z�ẵ�&��:�����{=���dK�m����-Q�;�p&����)��ؓ�$ �8ڍ����	���&Y(��m��ϕ��Y�r��oU2�OE��;P+��:rg� u@4���qԌث/���'�Y!�f|�تs����YB�H����43[�Mu尚��r8p�bDG�R��UM�N�k�ڜB��޼��
k�[=0���;��Y�@>�Yk���x�<jQ�ݍ�f��?��7ԡ�%�v�(L���.q�G;�`$S�
v '�ʄĭ��;Q^�&2!z!�s�j4�t{n� ϱ� s�U�l��_�P��A:�����fD��i��؜8_o�b5G�A�É��t�8��`<��XҌ	���}�C0��*D�ǜ��U�b��T���G���q0�v(������%38̡��Q{�f߉�~nw�o�6���xA���%i�7#ngpB��k4�����,嵆�-�տ�1?��I��N�͜�0b�_*@����R@ry-$?���3_�f������?a��15J�.<���MA�2m�`��S/Jo�����<���&I�7�V�:�T=��9�ʀآvn�/k����[�.4O�_��R�brфi=i�kT��U9CR4~x��~]�wI�|����<�ۅ�01� *�Q�/�t�d�^s\���ۍa���R@c�~!]��F�w�s�/X���e�mUb����Ϫw���bO{�����&�����֖��l������s߸���.Q�UdZ�k��ۙ/st�k���)gn��	p�Ҿ3:7ӥ��9��� &�&vR���jTUS����]����`��!�|v�����a2B`�@X�G�dƸ{̟q�Mq��N<��^�b���6��~doW�j:fY��� G��{�����o4��;�$�v�.�H�f7��Bx��xX�bW��^�Wb�3~��XLu%z} �-�H��Ո�J��z[�f�R
�{��u�op����k�k�McX,�N���j�]����f�i�I�x+E}eU K2��kI�E��r$���U����Fu���I�aԍ�}�u��݀(�3@<TG�Rݕ����@�])��9�v�D��N���M��]�Z'�'%o����|2x��/\w3�h�������/��[���=�����Ka#Wg{8߿�c9��
!"�W�	�ױ�єI�b�=bڠ���jHf�y�fe�R��ų������[<��J��cO3�%M�ܫ��'c�B5,��y\.ef�L~i���yq��{��
�$�߻���_��O����syp�����F�6���c�{f��<4��e�膄�~���D�#/��-&Ċ�x1`@������R�Zx5޸ar�e���ʇ&-A��XҊT%M�Eo�"���-ǟ`9x�]dO�JEg6��,uٴ.�v�D�[4cQ?� �ҽ��ͦg��Ù&sY"U�~�g��T����BG�Q��۬����������k[H����-
�������b�kY�w��YqI��c�@�N��}e��!���\��6?�����G߈���|��`�m�Jq8ԗK��j�t��N��I�;��}��gȐ��kr�;��Ƣ�5]4e��'�ߖ2�´��ͶG$� KR,0����8��TEYc�%����N]%��Mw7�2T�`�l�Rqy��j�7�I�� ��-{��^�zxA�3Su���oP.w;U�x搒� B�d����c�����<���6`�^q�F�=>m �����`��L4��@ �Q�[���g���}j9cM��X�U
�����`��U�~��VlG*��D���=�0��˞&��tS��G�~�:���pr!�Όu��Z)�� ;�@���v��5�0~v�<;@#j�c���UigZ=��FDX��
c��{bF�ϻ�l5���Fnv}��!d�66�v KlvXpL}��F�}�+��j���mS��v��S�@T���7ԧ:d9�RV�rS�����R�s��Z�̿u+��R����Y�B�<sW�F� 9N$h�c�ty������A^1�<*S|zp�_�L��Ѵg�d>��������ζD��r��i6>�*��~���K�?�R��t�ݳ�n���@[�`���թ+32��r=t�#�3^m�1�t�"�S�[9���?�`�Nb3��א�:ƚ��(a�ՙ;w��^CC2}�No�bFm;�+���U��o�C�\����^�}��?%�}e �X=�[ѡ6�o�v6��CyHCY3J��@A�5y����U &U�I��ʉ�z�Dn0������q#Ū�o-�������۔a��쎎I��N<��hq��f��
&/��@��еi[���S�F��8-ؙb�s�ݱ;��{*������&�e���[�[�"e�F��|�:_�X�mW{�v�eΊ֦�d�9�Z{ĝ^n�����18n���>��)�R}ܽ�-���-&^1�5ҋ�L\�}�\뤌���в*�?�k����UG���E���$��P#��/E֐D6%F��g��� e����������1�`8j�߽�?���+%[M��`B��O,�UN�X<��Y�@G [���_�����E����Ki¼����(��5����]�� S�ⵝb1�Zs����on��V���+��z#�5�t|FY"Z�����lri"Nt�&+���
S���h/& u���=Bg�@�$��£��2�&���`z���qݿ��H��N�8|�� � �m��SkѠj�G�Z�SJH�BڠHh>ge7������(�0�D�3�%}�y:��b��8<��i,�0��i�lSH�z,'�)��f8��E׵k4�wlvv�����IXG�Ľe�r>
*�������o���(��vt+�k�S��Vb�/��a����-�<L��T���T�h8/��R�7Q������
~��Vܬd��Л���� �Y�
�8���b>�4��!8�80�!�H�;�ۂp�Ծ��~��c������� )Op�o?`���k췢8	��Mdʟ*����C��`��Z��^H��pU#����W�дwk�˾c�����LU� S\���C�A���}+��a���M�̹;{+)+P��i{�)�LAN�3�8^�f�8Cpj�Psf���n��;k�̣��\.���)�����h9ʐ�gh-��j����@%�{@�K�/��&ڨ��q)+�����\R���v�M��zA����r����Lg~���'�)H�-��eTa�*���&�b��X��	���8���`;*c��?1��Q�e%;��	��"3u��)�p��|$�r���|���I<ۣ�P^��3�f���'':��Ypy<S| X�������y�{gSQ !�s���6ٓ�.BU�t��5t.1����ڪw�N�F��%�X� ō��|��w�����b�������RI%����Q����G[�G��%M"Z�F���!����yӈ^���s��&���������WT4�;	׵T24tx��6't���;��".�HE58�7�뵅�'w�j���0�4Ž��sL�7�S*�'HE�<w�}���x��f@֟n�Mk�U�WeAHg%��;��^�`��`P��]o�e��4��J�vw��~#xN¨��	�9s�0����c46�
}d�QG�����p�6f�"��R�x�\�-��Ob���ۨ�PQ�Lc��Q�}��=]F�����RCS�tխO_�����������0�C��!�T�.0��¤C�k���k�.�l��3=�^���3c�����7z	*�w#�[��RI�-���w���U�:/d��&[`D�+�<)�צ:��� �4E<��M�+�Ѥ/����qfw�i��3z/�Ed(���մ_G�z1I}@LU�.�rpĽ��z�&2S����<k��.���3:q�`I%�� �}�̿�{�@ i��7G��s����%����ɼ'du�ؗ�g[��D�i,�g�Q�{׀ш�&b�v8�V�ټMf�6��N5�>���^b;DG6��W�o��2��)W�� u�W�m��Y�Ase�K
L���g������� 7)Sy�h!�®G�ȴ�
��NV �uHE��}1y��:�4�`��<��nET������\�4�y《�ŁZ�-�����E0�7����x�s�o:V�C�8	����֦w���RC@?�5@8S�]���gF��K8�̀�Ί&]F���dN$Wx̖�����_O�Z�+zZ.1ʈt�TP28���?Զ�ࣗx�ڛy$���<�a,��io�X�~ ����C>A. @HOOwW�Ǉ�{D�
P���b������o��vpd���9�5r�'Wvd�5�"$ �<~L��l��#
D&��"��p�4z�'�^��#P�������!9I�u� B1�}0�:��8S�ܺ'� 1�2�b�^ I��7��,$ẵ|�NC�{�:>�G6na@��� >��+p�ԦX���)H����>���A�;��!1��6�씒�j�@zR����<-ǚ�ºpo��3B�'��R�e������tPf�oq�E{b�[SI�D������7�aA��3�3����m��le�#�e�X��l.���cya;�!��"�aE���+Dn��lC�g0����'����2m�7���-��yG�]wuz��J��[/�]f�>WE�喫���B<�H�k�ur|&��e}B�!��AvG]��k�s�j���Z�e&�g?�4�MBz��x�����7M�^�g�qb���5�������ὗL�[���S�k��0q!���T��{��TbW��c���wϊ��ϭ�"[�(�֩v�3�ɳ�~b�<�����Y^�,,��-�f������Fh���X3+W���?X���Ո������n�t���W$(�Am��	����&�"�V���},�648ˋ9�� �H)s*���nl��-�36C�t���t/0�
VG%r.瑻K�����[	9�츤�,��U�FՋ\9=ed��7 ���`��K�JMO�
G���\\ �Q���)aJ4�R$\�7@���/Ԝ�+��D��#�������@21��7?bzjbؕ��r�C�O��D�=M�D(����;j]gY_諭A�q�B+���0����m�Še6XI�gF�A� �����+O����o�:�̈́�=���0�-�w���^�u�0P�t���_|���=�#�H#�9*'"�dy�W��hfE��[�0�>	��C�ؗ��48ת�᪅�Rr�y�W��=3��ד�߯!��<`�"�f�[%�7��+W]�[#��u�M�Vvj�Y��ʏ
�B���g,�<o6ؿ�d+S�1Ҭ�t�/֖���_9]���7��A�M+�^u��=�m��0V�(&�#{3X��t�y%i�gvȣ�+ᨌ��o��R�f�0AW�7����h���������<.R�>4=�5#:1�ڞ|�QyŁ$r���p,@0��-�� D�HX���')����f�V�|5�i0; ���<�e6fC_c��Ǳ8t�o��M�=�l�Y(S��-�M2/����v���'\"w��bD�8rM�Bn��A{�5#�**FE��hO1�髊;���Xo��e�7����Z~dt��~ ?e�_"N�|ژ[;5�H�O^W�ڙȯ�F�%~�)��;��D���
��jd����n߁p�h)��|��N>��Ӹ=:A ��Wbݼ�� ��o�YL(��We~�b�e�ö9G�D����Q�ݝ[N ��O����Z��i��@b���mh`���q�Z�w�\�v��|�������y���e�%h�7��>���fF��5郯�b2ߡ��䎭�}��i����:ufI�����ь�34����7Y} �B�mD'�/�_���}�ƪwM�b��#����,K܎���3��D���#�2�C�9��n4PopR�ٽWN��Ғ ���U�۸-	y�A�>~��ee`��䛬7�� i��%�l�S��A��
��!����gJJ+l������
�L��5��N-!ƅ�&#��	�<m���%���oɁ�t�Q��N����j�{��\�$�G݂���~��L	���0�b�} ߶^�Y^�f���[(z�8����a�H�@ᙅ��l�_��1��}�ĵ"��|k�?2����^�դ5�}S^����4��M�u'�[�u��K�� ��\@��<'�_��%�+�S��c�b@qa��T���+d���oi}xb-�6�7�zR	e��g0�>��:\@�*~+�j(�M�l�G-pzXb�]҉���B �����֌>ZA�q�#�[�x�~�o�t�J,汣��K�K�s;x'V>�/�}�u�'���5�3\��A	�Ӷf!tDz4��W�;m��?!J�`��r0fs�5��b]G�b��[i���X��(}�o�Ȇ��-x-������!�X"��DE��bX��'c���>��tfZ+��K(�KoW� s�2;@[S��\`��K(�g2�j3�?I΋&h<��
F�v��j_(�l7�3J�\!��Q������Me���N���#"��r<.%����̨$�"�?Q�B[p|t5�>�[���{�V��+�T��=	g�U�S��Go�s}FQE�	�F���Od�N�w��x����3�CQ���oɾ(�,�:[M�ӹ.QH��^g~���U���G��z�f�T�l+���9��fj=�8����G8�y�K�'�H�}�+��O���������/�� ���rD�^	�`�h��VHǈ-�+o��b�O���Ǭ��p�����K/� 7	70�[�v[�(��tF�s�B%d��/�����ވC�ы~IV�X�4S��,9���J"��PJN��>�S:J��R\`gr��C�B�I����O�q�u�s�%���5��g�����,,G��w�u����&<��(DRb.8��C-g����Nli��̣�ϔ^�,�Ħ���HT҄�G��o�-��m�Ei�)	H�G�������MsT���/%X*��4s�����J�����49zrrT\�����W��3����7�DƁ�<ǰN���"V��9l
�mX�r���	�Ra(�`����=��M����O�k���VmIj�a�qǱñ�������K ��9�����4H�`����k��3��dyO��܆M*�l�x�}�)$&B�2W	�d��X�Q��z6���KS�7$��N0H�$N6��k��X��(�f�h�l���Y��i�}w�Ƭ������%󿱬���)!��
wwɏ������I0�(�(�s%z��P�2.Ci�3?����M
�xѹH�o5�ňT!ʐ7#5�֕b[B��������hH���E�ҫ�Hf���o·�x���evYU$:l��z ���#?qEv�y8�}y|$������t�@�@. !$�zƷ�r6L��E,��	=�4�$^x�j̙6C2( 1@z䜑��y����wt-6s��6�2e	�8?zoU	?r�Ûln�p}����+P.
��(�	�4'�W~������K�+.Sz�g~�?�+�E��s���D�Y��;ݑ3cGv6=�,��gM��v�!f���r�d
���F�A_���7{U o>56�����G]��`�zbQ��6|������d�2ۨ[��s�"Ѭf�� L-S��o=����A�|��[}g��\$f7��f+�,MI��8�b�l���:/��+풪���������C��o���y��%�?HY�E�`��7zdv��d�۟�����ԞָZ���D��Vj=���jޠ�x�ǫ�w��`�@��sX$;�v8&���D`;�I�:m��T�Y��Sg��a���~�r��a� І��k�D�[�����3v�8O�w���J8�!���V�r�C2r51���Pm��&\ϯ�����HxF�$��ݛ�� V�E̐�P�p��4��$�M:�� #����[�y�K'i5k�����:dAeJ�/�.���EE�33��c1@wLV�x�d�~T���d6����dw�0ܥ��E)b���ޢx�y��hi��5��fC'��e���`���A]���@5{{�inj÷�T��Q�Kט�M��9�T$�Ju�Φ�;�1��LbX0>2e���d�ό�}� [B�K����ol87Lp���Y?/ֆ�'w��[^���� k�p.���q��x���P(�0�PT����C�fQ#���V*��w7�xXb�_���^�j��ޮ��Ĩ�$2-h��-B�ʯ°��%庒�g^��k,�MGۿ��%=��@�5s�m hz0lob)����|p���b0;/q�5,8�����Y�?g%z��$���j��D������$�'4�a���쀰[ʆ����Z��x"�Q�{�f�4SCF�<맄DDtL]崙���g�Ð�:�Q��G36����o80�ˮ;��������ޠ(y�!|x˜�#��p_�g*be⊦_�j;�/��]l����D���h��J�P�k\Zt!4�Z�!4$�<�K	�!îhc�A�W`Fa����{����4%�"=����������'�>cEb�@���q�6�Z�ZXA����p��+�|�N1b�yN2�4�4�Z��Vp9?��1���&+�p� �������9cM�2�)XK�.{���˫�Pjw`��\xG��4K������dH(QB,<0)���?�#�!��k�n��|���c^�����E �hu���!��A����X�M�Li��O�I�~����{dG���+�˾X�IeÕ[���3%����4Y�o��kej�r��2/�d�wC\i1ӏ_��=aA�:�=U����)�GP�4�Q�-��?�^���F��{�zg�L)�I4[����k���T�-�/g`ȺX~�0��P���t�@.��ݏ���f1T`���3�Y��g�k�ɉ��G<���&�Q*������V.�F���^],F��kk=t��uT_�0?�ү�P̡$�q��!�(*k�62r���7D+r�,h����MCCXӌ�7�IX��hB'><W��%��L����Ķk�@�]k�{9�痫3}p0V3�+�\x�U�R���!�TW�u��r�X���N�6{��OL;U�ʇ���`p;���}Ż�/^v~���Rv>����yl/T����_�ܷFk����	-`k������2�~�~���sU㏀	��#�)]��{�"���QL���d#"�8!�
��zp��d���r>��D�����{�Sm�ɩ'.c����"Ts��� ��	�|Z.E���Cs�f�+vqo�܋��o�)Z�;�/Vf���y\A;��iB��4ټ]�|))����=�ё6;�/�S�gzzT������D{���x����礅O9�ɡ����� ~w�5��y��:��)�M�q����ni��>�eY��	��Hh81ש���RO���X�I��|/�j�,�a-�;�,P�i�C�Ձ9D�����.��l��.L���"�qN�E�px\��IqT_&���4?	Bah��h�a��Z�RYlfؗ��\��Ƿ���M�4׎O�kb47r8���a��N�-މ�jRQ��%��II���Z�9�Yy�ޓ_T17�H�iDcY��팑�)m��~����B�t||1��/�k���AMp*G��3-&���c|k�AW�a�dR`w�?��)��y�y[Q��s��vI�ϣ�$[t���8���:^mQ��J�S�[��ƪ�S�f?�-J5���.ɠ�S7I��#R�¯��B�q�T���g�_Љ�/�vlk�6��w_��Ƌ�SQ�hAZ}�͈V�)��ט]�B�i"/x�Y��I�b�F4M�Hd�e�OB7P�Û-}wI$E��yB���ٖ��A�;�I��5]L�2}�nu'n�_����asBG��P=�$c��o�\U�� A�C%�C�A!��so
�I���s/� �^�f�'JH����'��ܽ#�;T����}���@=f�\�`n��FJ�����B��r�,�@���,�D�8.�Fe��J�B��H�0;Q2೶�� yhxP�(��mT�``
�`��#�� YJ���B��aXQ���際	�gQ�zT��c&���,��c�e��ǿ��愖Z��������w&��N� �%��ߴ.��c�����Q�s���7%w�&>$�J�(�9?n��T¹��ǈ����|,2x;��搵�|���'�n>N�Tl^��(G-u�azd��Vr��y�#[��VK�/3&��3�ʫ6-P�?�R���L���}g�v���7YLX�L�EHn��!��U����H�d���NE8uH?�3�m�>)���_�K�L(0*]GU�I[���o�ݡA�ߊ�Rpz��â�rxi�Ե��3b����%�r5��m"���p9�d���{�W���"�j&��2rQB�"o�MпSN����7ǵ��-�Nh��~�F$_�f�#��G/W�e	>���ܵ�T�����B��yF��&���銑UR{�&j���Ⱉ(Ns��Ƈ���
�$숱]��U$��X�?p|Q�c�hn����?���;�b�m��i�2��tqI�X�jW�]hc20\���$IB͍����H��jT�a8x�8,=�e�(Mm�da�{w�S �`��6�5z5Y40�{��	����R��Oy��`:�btV&�#u9vF'h���f��h!:Թ;��6
���P��,y�yzZn\�4<���_�ۘ�4̌�x���Ό\�?�w$�[D�ED�^���$j�|��s���n%$�w��i��^�G���F/��(�E�M�1�)����˗]�I�=/	U�c�׬��X�u�2 5�rV��K��L�0���q�YaJ���n�e��)��<wff_�D{eTm%2���&A���d���2�Kp��w��ap��������s�OK=Oխ{�����/�
h�Zw�."��n�3����NR�.�Ү*�{x�0v}Zp�3�"6wc`^Y�����7��Њ��v�r��^M����l��(���>���]��'��ƛ2�D_O�g/�GǊ΄A׿�啜n|��-��GU�:8i��J;R�8�˚.�@eF���
ktÐj?	�W����])Q�BNZȮG3���~s��͉$��ԏ8�Us�̶J�ypQ���?KhQ�}�&߄��U &<<>��}xU��-5�+Q�G�Y���FH�R]]�����R����t��.�H��ȁ��E�$�9~�u�&N�8G���+v&d����?f��u�tD�"X�����'��Ip�>�4�[j��K�I�9PFz�w\�j�>I�lZX�T>��O?,U��\��O���H0��c�*��E�{X�ό�;B�).�������m化�|Ae������;��l#5ba4]
ˠ�v�X�TTP�k✔��;`y	-��Mݼ�C}�u����__��������%�4/�T����9}Ȑ� x�6��<8��>D��৷�kX��A��`D��ܓ̖��̲�u�L��9kY2����H�V�ˋ��5`a_�6�*;��K���cq
�����l��;}�-�4
�<����ť���.O�ք��#��������Ǘ,��G����&��V-�y��k����?ZB�bN{f=k���ie�_�.>�O˺��
$$+��V��r�=�,�3�f���H43���s�c�y���}a����ٴ��$1�k��7�&����ÕP����C��M�B�sQf/A�~��_/s��.IJ{BW����GK�"T>�1���$o*�1Ƴ��QQ�!�y55p���d]?@�J�_}�	����Zlq�P\��~m�%gx?��M�
L�"��T��#a��Sv޿�@@P���V�U�j��pg2�KL^�+���{��}�NUC'���{ל�7k��'�L�����VE�6��ӊ&��o��9���S���W���j��ִ/L��LAB={�YO�[d[8�[�w�V+)��J�=�=~��Ȫ��x�;����b:]/��/Ml���r���S _zF�bzpx�G��bT�0� ٠�Ð?;��5��ɩݤ���Ȓ�Fh`6�L��X�[?��C�������ԧ:�s;zSg��*�o���O�$��_-y�Ϋ�J���S#R+'!0�����H����X��}��M��˚x�~}��HN������\�ӂ,�:�W�H�#��us:+�8��f���4PgQ�vNL�4+�Z��K@0M>�x���z�D�$������D�Z��?��_0)�gZ���3,CpX�ݯQ��5��,To=*�K�/L@��Z�S��l���������<�2+���L�r��s����M�Kh��D�
O������R�*&bk'ꝅ�+��o�ޫ���
��r������Fzdj����̑E��;�\��Xi�ŨiM�og��5���I��R�&Jdw�m8��l����P} AW���*�	�������HkxX'��|X����9��NV�9ZĎ��d�
q�.vgrգ�L+v"lȒ�6�����3�+mلQ��Icf�m�G�Ǉ�S�dY����(W`!i����/|���³Mq>M~0��+��j�D�\C���B�SY�W���{L}^p�^a�	'�u���2汲�晀���R��&����C����I�gzmm�л��/;.b�P�u��T�ԙ��e�if���ūi���ɇ?F���-�Գ\�<���I`��__f��ã
�����>G�\�^�¼Q���y0�RQ3��Z�q�F҃W��ͯ5�v�V��2B{R����+'`#k]ي5���fc��.f�V�/90h��:Iq$���\F:�F8NW�ݓN��Q����2�xx�(�A@�ڞN5e���}��=~֙,��s��}8ޑY�=	����FPd�IVDE����/�)HrX}��Q�\Y{���R3R���hWeRMb��Pфw�""mۜ��HEM�	���C�^�D�<�rG�$1~�BZ�]�y�ww5�.0;������jc�:�?�4��7��1	�<'&��XLl���=2���M
����K/���v|��<����2%�?�
�[���Q~��T�8$�a��L�;�߽�����Sx�|Ͼ�����rF�&��d"�"��ak�1�X7�l_�yF}A���G� �A��߳��MT'$��ѡ�P�P5N�Ȕ��"�	sɨ��>����;� f|���$UlD���L�ë���{��i��z-3*M�f��?��}�up�'0�-��[J�tP�Y�>>��R%{<�]�ɫ�:�iu�u%��f�eu�&�2��1h�g�����G��J�/N|�����bU�{aԱR/�}�&�r�lSV���*�ei�?��#nP�Zb˘r�8���m-x% 4=��u�f�'�
N��;��?�. �rh�w!;(���] �𒔙�i!N�K�(-"s��x�vF�\�W���s%�����7��)�5QMh�#��G�M�3~h�]�9Q�E�"V2�4	Jѵ��U�x��R�tQ �4��������C���	0��?lJ���+,D�Ҩ
�Um��0P�@��Gm�+.��1��<��9
gR�_Hc�,G1���T�J~�q��FI�%jT�-������ժ�	�!H�)��5���(�6C2�<S�ヶ�@�鼴��K�����|���Z��~�I{c��&�-S�*��{�n���>G���BKU߷g��SVO�â�3���~�f��1�#�W~r9�?�,���)F#���A ����(�D��6@c ��x��HՑ��^r�bkә.��Iw̡�m0�hPo+B
�U�Wl�b�w�J�͡��45��#*4�q��q2� w�.G�DH�>4�=�Y�ť�(���0�4Q�V�����@s׹\��fu	6�Q��%,狡䢰21�W~���f�v��9��vA�j�X�I&�~铰ݔ��08��g�:��&}�}�It��0X��S<z2Z��[�ϝ�I��$�7������o%�����ϧ�W?�Kh��B1�&�C�,wZ�/�-�mC�k�y@��_�h!3���]�T��Vc��a�D4^Zd�M�ޑ�:���U,����)�k^S������uQ+�G�*4��t{�i��k3�l,d;+��c��׏���P��B�ϧ�VEg]�3�f�u�^��B�(3&���;}jm�<��x��
J7j|UaI�5&-bL�6���>�����^Z��X<\�;T���ɿ�ӎf��L����9���;}�81��:�@�(�p5��qY��Ӵ�!уXǽ��莦A$�N��#RF��Y�i��u:j��M���~�x4)���抑�\S������(�PE�ҽ�'��%M���¥����঳���#`�^�{�G_����z�4�uY�}#���X_}/��ZC��R�@����ғee:j��N���$�ϙH��$��AQ8D�/q���G��T��z�K��U>oaZ1`=8_��i�C�f�ƁSϻpt:�t�n��3��u?k@�<��M�
=�\T�Ól�bi�^}/K8��dYd��Pt7=9؞�A#ʄ��t� �#���Ѓ�5�W���զ����܇��r�I>Ofg�c�v]���nB� �e�Uכ�Z�}�6*��"Aάqa5�"!�����|�V�C*��ݢ�'�e2���op70ƈy]�g� ��JC>��{�|��N3E_����O���vLH<�����-�VT��w�g;���Z��%�yM��Wo�"j�ԕ�G����XH �A�Đ���B��Kp�D�tx'}�M����գ�����<������g�]f��㡼EGe���^�l��׈z#c/����G-��q�&��$�f#ަ�%��B����󒉌��[�20 �mʅ>������Us����b S�T�}&�I��z�I�����Q�bCm�I���i I2z;�q��7($�8�O>߸�5�K�ϲ�n�f��h=1r�ʭ��|����#*�#uP�jΡ�5Suf�-��-��lmeJſv�b ^�.}��="��p��_���$����j+2M��,k;*��o��pS{_j�Bȁ��ҍ}���n*���r 9%�.��q��n���05�_�0����a☎,f���������77�G���^~��>9| �����z@�]a^i4V�2�=xύ9E��a+,��y�DPQ"�nɣP�ᜫN�g3�7���ld�bx��gW��-;N`�><��s8�\9���֌�V�v"�n�X�"�K(a�F�?�a E�IQ��ןܡ��5��	�:Bb����>��:>6ԅ�_@2�����d�e������w�
Ŀf��l�x�EoE�:K���ʺ�,�_b]�Vl��H�e|�$����;���{�..��.�i�a�:6j���F��ëW��:�n>��)��[e�X̘
�8-���Y��a�޻�_51AI��3��A�Q�7/��%����l�6a��/F�&�룔��U�t9�f��Q�n�s6���3g�N�dކ7�W��ue�i�M�Lc>��T
��ѥ3*����率n�O'AKE��=�Lݤ��d�t���@pKPv��%�=3,:�Z��ɋbh�����WIy����6/t)�ᣊy%�>�T���(�{	����΃�8:�ru��ۚ��akN�k-[���[�eik���s߉"4�����8~���U��C�$�_(���h���K�10��,�H+z���Đ��H�*A��N�#ְz��������w�`鸠���|D)P>}�4��[��+�	`=�)����$��+�o~kZc�P���Ľ�2�/��,'pph�(�n���T��AX#.�B�B��$q#��N�z'{���h�oe	�aF&|Q`����#F�{̱3����Wه�$�`=��,�h!�=��h��?b�/T��"�HVYxT�<��Xd[�_������x�b��Ǉ�4Q?�����y2U�t؇�-�r�Y	�I����;NEϫ�'��2[�H�q?���#��P�!��_�:%��Կ�Q�ÝcQ����M|`u͐n_!e�I>8��߳K���U^�]# ߖ�b����UT�X��V�W��?&��	{�v8�1��
��ۀ�� �0>�P^�X%w������V� ���'簪_���ݏQȄu��$GH�ߔ�.��J��|v{xK��ߜ�85���,v>���5~1܉_��f����t(I�dq�Tή�I�`�^����)ﭏڗ���_�:�!a��y͡SՉ�58��u�?�v	�3��5-�ZF�T��.%��_Enj�0-��R_�;U
���\�qE�ȟg���:���&�P�s�ț�������Oh�E�h� �nW����{���6Q�M���ò�l��h9����r��C��Ѻq���H �s��jƴc��Y�vxx�%�Ċ�0:��Ǳ(:�|* x~�)�yi7��L�އ�����gٮ�2��X���XM�t��o��Q�v$�]`�J�����o�z�XOJ�X*m�1<oe�D�I[�42y:G��w���3���L;�N�A��;��#g�O���WKy�~��d����l#{����%_����U�G$�3��?+@��D��� ������{2��ݤ��tܑ�+['�Sp�4ew�W���N^�S����z��a���`����>��Ǫa���MA<0�+7��)����*�⡩���������6�R\�!�Q֗M2�C�q��w=ר1�b̊���G\��!x��#�z�O�L�T(�M�gh����C������ �-�^�3��;p|�
5ܓ����� ��Ԋ��bH��3Y9ހ����10�0�+*��� �n�S`��H_����i����1�79|�{{mpJ8cO�ar|�6uN��~���� �g�>!�2y�yy��ΰ��Ma ]���?��%���j���'zS�2����J����#��b*|��h�?�+�4�y��[���V9�G��>�ќVn���D)`�s>4NJh��m��z\R!��ΐ���zo�@�%��f,]�7�L�;��!�_�b!%����-�_Z_�u"��7�����4#&���έ�G�����r��a�v5t|g��4T��;VQ'�E't��V��w���J� ?T�s������r��[2�$#�p\5�$פT;#����& )Q��0�5`^Q.5�m� M9$��l�G�����~e�AS��Η���Z�s���?�[&���Bz,��/�r�� e-M��s�<�hX��wsV�����ɥ5'����(��_ �H����M��+A�%^n��-���Q!��4x@=K��|� �/P��XG��(G����� ��xߙ*?t$_rL^��(D���T�,
^M�-E�_ΣBՉ��BU!I
��{�q}c�e��A>h������l1`#�碦-��G�e�rAV�h:�G���Gd��ԇ���Q��I^u�:��.d�|���]Ҏ���� ��������.���������@�|���H��&�T+�H�tR�]FR}O����f�}��WϦ��_���Y@O6�f�ERt��_~�z���xo�su���]�ʯ���� I� �2��m�C�lI#5������sR�v
�Xt���6h�����%ٮJC@�_)6H"	;J<��*'�=��F��H�-� E8؃t����#��5g���� $|�r;̮��V��d����ԥ�-i����8""?���ӧ��t��a٩%A*%�UV��㽼*�>��?߷>��W�Y��n8o����0��Ώ�T|�oA4�ᛑﲯ�Co��i��/�m�rq�? � w9 �M��\�u���t���obq��y@����<�[����|�{C���i����U��h��&�&0�$%�7C֫�=�Zj�nGؗ��W8D��*1n��	h�ػ�/vi��s�
�;���-B�ߡ$���LQ��rπ�p}��K��h3��?En���iꋙ�_?'����1�MM�^�ĕ������OƇa/5CYA���oj�?�8vy�<��#:�}�$���h9;`I���ϰa�8���
�	���Y~!嶆*�ŵ��.�_���G��!�%e�(#��lUJn3&0�T�>���N��>M�*���;��_1kt���$�KC4���S_[��ڵf]����抌Js���R�#����Ֆ+^��EB�e�gv��9��x�2��,�`ѿ�y��ɱ��b"s��ןu�7 ��G=���$θf<$�">n����V~�pHg@7WhG�E����!�h��+�R���<�<��B�'D"������?�Zi)������	���,��O�=�HR!Jiɐ����n�����G�I\�/���h��#yD�F��p Ѡ*�i�������m��KK��!Y0 ���Y��P�|��Zi$��逘1�c�}~�J|��#	`6�֣+��V�=cq��5�� ����O�.�|��{�Ӹ��G�K��6H�|ǭ�~ I)�����=�s�:C86#�� ���^�<����/Hط��;�N��b<P]�RS�Ѕ��P
�Ʃ:�9�5t���CJK�*�`��u֗cޥ�#3D�(����oI��{��W{U�h*���q�[��S��5�/��GhD��h��C���(I٘ŷu%��\�cԴtd�K&� Tw�ʂ���ټ	�Q�\~��OF��
9��Q�uq����.0l�H�n��un.C�ϕ�L��@fC]��=l�X��GF�m�Ϗ��WPu�i�U�@N@�$u�I�wB6{JL�,U����}H0,B,����)���-�[����ˇ��Ʃ"p�`ع�_8p����8�3�ɞ�7z��{F��UL�����ߊl"LB���_f��8����nE\��g �Q�����b���`\�����~ t!o��ީ贐ԫJ� A>B�C���L����qa�{�PJ�rfhu� 	B�ax�Q3N��c�إI]w��Gj1ڥ��W�#�"�RdL�G\r~[^Cڴ�*�@iʈ{�I������E�?Am�+�w��;�G�C�;�h���C����J�Fp�wP�C�*��Ϩ��X'���������cǻ�0]�������v`���̌HB����qs�SԻ���S�2t�P��<zp�9�쩧�Y	�W~KE\�S�L NI�B !f,D��Tm�?�pيF%Zd�P73 �h@�*.��w�a���.꡸�)ө1!�^vȫ��]���J���!Y~:�]��,��D���A���g����Zmw)V6M�M�'�P���!�]�P�S�� t����%E|w����6�}�`v&�V����V"�~%LT�IU��(��A�f�=k���;=1Ċ'��HS#�`.���Pr�P�����ᰕ��~�)�*�yOA��7qҭ�՞�<:��d!�W��4�G?4#�I#�V����nW���gDk������D�'����[:[�#���B��d�h�Hyh�C�j��w�Ȧ|�W�1���^�)����Bo����?�����A�P{q�������B-2�����v�y{F|;M�&��b
��Cn��(���͵5TPf:�<�/��.��c�3�t�nZǵ��BE4��;5�^��G��][h9��Ob&����y���Ub�!�dbeA�=uWM9?P��#���~�r����n8#މ����b�\�C���7O��'��E�0�Cqe%�y=�xj�0�h���^�BO�	�dYY|l4�C���v�n�I]	�H�VY�ut�*�ћ�T�n@]0��0SNfg�|���,H�)�ʧ�0*�|J����xC˙��A�( kҏ�X�z��l���@�a���jY���?d���w�y��{�Gq"�x��ҹ�:�������?k�o9���`>n�^;y��g�M��	�~��� 	��˲SZ�� �k���s���W��������B*r=K<;.�0&��
z�����C O%�,�x���]q�l�`Y�\��7���;[����IǏ ��t���i:f�z�#<6�FIvBxE�x���j*��_�Y�L���aEg��)�o&t/��b������mqwE�|P��	MPW}=�G�Dj����->���K��N��?�����Y>a!c�;'W,�y��.b94�}�ڿ�6�.»w2}ח�y?h�7��GP�����JY�/ -��jB@��Ӹ�+^�'A�]���X�"�j�y�0�����\<.�-7Xjlj1h%U],�����&�*C^�ۙI�7u���u;,��p�}�R��������,+cˏ�Yӎ<=��Z�ų.�+[G�xB!��_8H���'<�j7���=�Ϥ
�P�x��2c���y����W ���`t�ZzU��W��ݯ����m��B�������S�3����q;3�\����,���Mg_i���Mg�an�������*Nwj"��P	���FbbIZ�S�W��T�]�l��?U�'��˭m��:�p'�ȵ��>��%��a�`���ވ��vF��QdO]��ɭUH���$Y�?�I�a`���MU��n�����βFH����	��ط2��ܦz[�
�>)q'S�{����q_����lф�/2{ͲR����fFH/�	�ozI�r0y��p�e�X4��H�� �X0�<D�����ܹ[���[�������w��l����{�����|H�^^�d.�no�GR��)�pFp�1��Ь7~5p/�"��S��vd�s�D�7��7#��$��H���Z��a��6��1}�? ��� \���ö����$^�!�j\���⚥�Y�/5		��_���p��y�piNZ�!�5�1������[2 	��7 3s)�$������@~�����2�Ŋ��S=��{r���tѓ^����{9��}m;r���-�m�D;n�����l�4搫8���E���zs����l ��#��譼&��
���&cD�îyb]l͂��[�B��El=E�V�ӎ������a�=���ߥ����$������sP0(P�{���}�El�U���s/�Qd���nX� `��)d�=��J�~U���o�F�<k�Q�]���.�	�A���O.4q����d"��6�q���E�Č��[�l�� i?��1i!�ә�Jc�9�g�t���jDǉ!��ڋ|bz�1ڵz|��-2�8�(���x�Z������ot��&:0�{4��:�_���Ɉ�r�0#>�;dƦ��L���w��'ٮ[�o{B����˛l��7�z7�`������&����a����Ez��J
||ɖ&�v"���,�U�;lo�p��U,���/�g.<���"�0$�		A��O�)�gX�7Vk�@V��f����7��Ƿ��c���Ϭ�D#�Be�͢1�r�EyS��l7�q�|��0x �5�c��-�˟�{�{�,��.v���Y"�;��(C�b��I �e���9��,�߲7�*[A�ܡ��נ���!p%�,x��z�e{{�"���A��zjӮZ�~�Z]���봞��r|�+EA/*F�W��E��g���t�Y�V��C+{7�v(�q�2��V�PȆ�耴���f��zقl;�H݆��d�nT��O�^=���[ڷ�°(b��<1V;O�'��175q����{v��_������c`�_ u�l�L����S\��-�ߨ^هg�z�+�v�U=׌�
�5zU)�l@ ��qR2;1�R�lVxR����h��H�WnN-�NkB.O�5�iB�F���۞ �4c���M����u��5�M4V�n�]���Ր�!IZ�x���*`����P&��U𪋞�[jjw�H��UA[p��d9Z�E��}���B��I��F{8�������6=��^�v޵R�E(�VݽmN:�s	�9��q����o��h����k�k��������/-X-z��#"/;}���J0�J����`����Bb ���
'P�W��C%��tV��������S�J�|e���T�ý���~w^�o����F0�m�3r������q$H����&'��RV����t�<�y���,�j6�u.�I�|��.c����k)ͨ2�*�݉�Io�sډ�ӓ �f��CO�N��$�0>m$6������M�Q4!��y�m�e�&��f��
�=�]�W�agW��d���.�W�'[�p(�mosA[q(�T/�;���3*-�\l�A��eH�6��V�2�9�x�n�X��a���_���s׸\l�uӇn�@"ԅ�8f�U.2��KN��	$c�쾣���4����U�9ў�Wm���a+�B(��c]�5z�n���2���Fy���w�����=G��
,��2�~�ۗ��ᪿƀ��f��m��MDL�C�f�����=)%><c�Hͣ;eӽ�>ND��*�����d�m�Ì=�J1'����`�V�t\i[�������p %[��~��1�k.�1h��~ʓ�%�<���=˘?N���*���lC�S\�
?{�����=�ώ$�����'�!��oΏ���˨iϴ�krvPd5p��P�h��IR	��m�9Wց1VE���++q�ː��߃�&/#����74���>�W��Q�K�FD��?�����#:��m��MHb������x��GH��f�BS��$���-R>�(��Q4��g�]h
�|�X��0���23��ܢ�T�d��r�G<Z/D�Q�7��:b��<�YX��Y􆥠�LVL`�1���K��m�����#�s��T���,�0�n`\\n��o+)������'�T�>��$Dju�7��_4D.Os����d]ԊAK����m��-����i�aH�~_���l�ھ�P�Y?IT[<���<A����=��.��@��F�e�8���M�G���j���g�^
L��3ʃz����<]JG0u������*jC4O	kT���jH�_eu��OPB��"��\+�������>q������2T��{
�q���x�_�L�.c��
��/���V�b�����ӥu�H��l��Gj�Gx�\#��:�ᶓ;	��2s�%K�i�X(�'��ٿR�BޞW�C}���:b�1fH�!�sb��a�z�������A�L������ݭ��?���͞�н��e8��(�e�ߡG����ЛC�����n�����[id`�h��lݾd���6O���k� �l�L�C�Z���GM�p�>o6�M��ѱ��"Y��YNl;�,�q7L-�u︷�4��?{F�F�@/����Iz�f9��s�u��H-�y��*i<�8VF��1��'VmC�Q6��{��/��n♹�����čo��AR�{������.FT�:M'�o�,��ҹ��{��;g��b=��R��)�!%�	-�kd чf�#���')��"�����+�z|j�I+��!�����'��v�Ϊ*�-^��Ѝ�C��^�~�A���e:�n��@�J��l�-թɪ��1q�6iges��N�g1���]�/��l���܆�Q@;�4��}J���
D*_�7�.$�υ�K�*d"_Aݞ��^��+^���2���V�Ĵٸ���S��ռ�͢��!{7��74�]��.�:`�#��{< l�t��so>}cO���GNP��KQL<�w<<�gVu�R��h��,]�q�>�0���8${T��٧Gs&WB�N�#��m ��`�
N��k���0���}����6��vk�"��[�c�����~�m}��?;2]0�A�K���᧭7������l?�2"~D�e�O/��(Jt0�N3���G�vf�M�!�D�Y���8��/�]'ʃk��
Kc{�xK� �J�dd��\w^��U���k�wZ#ވY>�8?�WD;�|	�&(��߬g�tЗ+�y�ڧB<�w����(�Dg��g���t�D�<.4�|�Rv�?7�Q ���Tm�1�|�ۀ>B��K��H=�n:����<[�'��F+�T˛d��b� �ͮgJv���]d�7�%p뱞�/�(���>�Q0�Y��~�F���h�կnq��%0��Ԙ�|���eE�U�A��ׁe���%������5V��i?)p���F����s�YBS���~�\?˟�$�i�n�y�EͰ�\�y���eTxpω��7��,��mB �#�;��i�D ���-�����E���M��(>ͿRG�z�u��lgD�������|�4��%M��/�=�q�<g�)�xӆ��hK�>q֝�)c��>7�j�sy.W��k�{.fD��L�[=��edG���3�'��#��v�/y$@h��ѡ���,+��A��y�Y���"�d��}������Yw��PnƩm�z�#�T����V��q3��<Өw\ϣy5Vv��M���E�%�t4>�j�+�<B[r��ONo88�Oc�AF�4�:cM8���P|{�7݊�G����[�x^%�+JM��`[%|X�w�)��ͫ��)q��%㠘;-A~P,����[U_��C1-�Rva��"��d//$1ρܸ�L�KP`���)�Z��y5���z������C ���_f�疈��~�P�� �｡��C��pb���jPN}\���zBH�#�[�Z��w�1�aVoP�xZC ����	�eƗŮ�"Yze��1x��ޱD2�l�5@n竈��|������/K��ZlU��k���Y�_���4��o,�ۏy}{�co��f��q����n�I���!5K�O�#�Lb�b�c4��*3��!�Y���[E:M�t7�ם"Y�Z�.���$��6��?
P�t/���2���ȿ�]�z7OU
H�g�-�4���r�-��69'16��q��K��/f�'�W���ݒ��@י!�Zy0^0�9�3����Wg��(�Y֐�96���g�uU����Ųj ���à4����$P��O
�*F�����;�s��j
�J�r�8h��}i!z;�E7�����!&g��k	�K+MN=�l`�Hm�قv��~z�Ѐ��/�Z�W�!r�>O��Nյ��w�w ����0�f�HF*��S�m��7�,�p��6�;�Zŏf�J~�"g^󸾇(�������Mԕ���w��<��Ǒ��e���d�v����%�N�1Ӿ�}QC�P��n�7φ _F�E�"�@@^��+,�%�K�7 ʫ�'���L.�+<I�t�A��(h$��h�S�^:�|0�#���PR��tF.���$j���ﴲ1g��=jq��\��I9q�P2��%�B���Q������?`�(�
��9�_V}��w 9�G���K��IC?�]�2���J��ު6�M> A����#ɠ�h�����C���%+��;?נ���+<?��;n!W��g��PV����4o%ݠ���x�VE�v��w������WH�&H�D���#�@�:Rh�&w�"�����H�?���`*�!��mǫgq[��\�Ͼ���^��a�xTE��Кg��D�|,}+҈���b(�5�A�k�p%�殄5��X��(Wl}�Y���"�����Ǽs,L�Hig	�,�v��0d�k�?Ʒe�Vv�@#�}ǰ-9Q��t�h)������uH�r ΰRw��ɥ�֒����7��eV�޽MEޞlB����قt4�u�mh�R�C�v���'����\��
�AsU���([���g�	��������u����<b.�Q�p�	�A(o�$���Nֲ���M��+���T%FY�=o�ugaഓ�6-P�O�����q����o�ＣU1`�.U���qɿ.�Ib�½�j� SDv�2�m��3�����C�\Q@�Cē���_.U�}h�~��,˨(���Ν��Y����Zfc
%;3��[�@EgB���
"..~�1���QUh,�?)P�����	(��;$�90��]2�GP�)\��h骪�v~�I"�kE�I��
� V*��&�TU?��iQ�~
	;�7W��U��|��@A���΋� c?��x L3�kZ��}�M�34,��E���)	�����u��+��{�D��^Zo����ʑ��wE���\�E�����uV�����M���*	�)gzs���_|�R��b�����mb���B� �Y�V�A�E���<c>b�	�(ɢajԣ�B������#O�BũЃ �b��1�\'�Ob_}�>C�]��S�l�b]�{, �����A&�{f"���5��w�<�ӂ"�,�;*9v�!l���[���k�>��$^�"y��t����* v�?/���x��/H����7�A�6�8Eݮ�lA�������w)VPҠ�"�8�I��r�4�k�X\2��ė�X�)|��ĎN}d��;��4���o���,���xN�H��OnK����0�̍{])a����~w��8�(��f����R�$o�JJ2�}�o�kЎ��z�sOk ����&ms>�����v)�q���,?���Lj�pC�,��P&PD:y=�GH����>�8Қ��A�΃h�mD���Maz��"�"�ޞ;��:���X�ح�7��!ȩ�ﮜO7`��C�~���K��Ǳ}���#���Rs������$b��V�1MY�<A!5ɅU���Oy]����*�r!^�)�d-@��V�i5x����("��@�hj^���P.���9RR\f !�N?�����$��ϳ�H�[}S!�e�M2���1[cξ���[�䊨<�G{��p���#����qB[��	JQc_u쌡�<8��s���
ԕh����nG�;>s;�Oo)z�-�%S�/������p|�R����B�b*�*lZs��c��`�-��D���P�Zi�X���|ՙJ���NB��??GM�mH@�Ch��P�	b\�vK?�K���72,�Hu1�\�2�%Xl߁�Ps���ҿfaH�Z��G,9Z؍�ДЬI����8�E�«��k
a��Qg(�k�Q���f�l��vbh��~7�9z9w̎V���wT��(R�gx#կ�My���w7� ����F��Rj�X���X�#n���Q48�X����	Ƈ�,6�l����2��?��
E,�OUX� H_�R��#FHoqIIw�\YMM#���{��/Ah��~l�kh�v�2*�.a�)��.���Ejh�@@�[���@�P:��fhAR�o�=�;�}�Z����[���3�~�����ޛ
�a_>�yT���%�D�PІWk�����D��.&�������ӱԬ~6S���?ƜJ�U�������<�o��*e}�S���,���pmը�T���ܦ�5L�}�^����c��{��ʃ�"�O�Q�LH�xC	MD�U"��rld�&* �z"�������v��bnL�B�#��7%b�O��I�B��Q�y+՝�򬗒�X�	(���N~����XE�r�	�	3奶����{7}o��~�_l����U.���<`���"�޽MɎ���X�,_�R�p�6.�E�2E�s��454n���:�����w���C�F,eGU9d}�Pi��1��zG�0@���a�Qj��u(]~}Κ��:2!<�����+���ۋ�P$<�n l���m��,��,�� j�l�2���(γ� n6��(Ty��\��J����J��M��r�=��JpI�'�NF.$�QC����lx�20x���>?��������9��λ��vp�[^���cB�'s��m����,�P9�9R�b_캯L�Cs����4���TC�$�Z���~|]��n5r���s���_�,b�wr�k{�b��>`HB� T� ��i��4K�����K�ÿ�_kt9o�xv,ui��C���.�CX�Y(�L_�(?~U ���e��;kS�7W�5Uv-�w�{�E���b��}����o�aO<��.��=e{�7:�\z���9E�69�0�N0䭶S�^�:^v�&�~�A̸��j{�����������J�����rm��[�_|��®���9!�����1Y(�7�Y��O������g^��ݜ.��|�ظ@�uN����m0ʠӧ���j���k���p����\�s�:��5��1, ������􄑛�A��j3������fw��'��X�3���� Ez<Ѧ��f����Ĝa���k��ޱ��_����q�D�Y����֎/��Z��Ǜ�}|^/��n~�U���;Ǻy�Z��7{<���g(f}^KrN�2D�(��S���_W��%48�;[�?���<�!�3�&o=D��H�؍��@��M�Ak�����b
N�M���o����e%NL4N��J�]B�]P̈;�x}%hI��c	oY�?���5Һ��<���>����)h�C���q�B`��DA�qO�C|�e��?q(Eq�4�a���y����VZ�)��+2)K�]�����MISӫ:����K����(�����ؾH�]�Q��E�z&0k䓥,X#��-�w�V˘8�A�"�(NePqm�^9�87h��]6��n��N�܎���h�E�P�c�i*C����ֱ��p�!}J��*$�_�S���fg!�����%��M⡟HX&yG�f�`,���MTa�O`=���B�6I�*����lh��S
V��g��ڵ_o�/�y �Oj�5c���2$�L�xu�K�z�z\7��Ժ��R,��2���x��,����J�՛�3��񯨇����g(����y�c�f����r2� hpT�TUp�~�΅�R��gT��	�T�6��
��˃yE2�d�x�.�	�O;i�	b��n��K�`�\�X��bkt~y��!u����[�fB+AH\�:�����͔�ep��	>_C�^줏e���ͣf��9���)	K��O]j�nH�E���CŖ�����p�f�^˪��~V��qH�](1�N�I;��Z�9��y�EA�>xJD�������4
�� ��*Nڌ���I�Y���)e}n��Z-���� E�H�&I��+g\8���n�a�2�� �� Q�A��T�F��)�N*/J�/��V���(�q�:�c�����<n����e>J��gc��t�,�C�]�HO64/nV�u��g5�Ѡ���ĵ�Ej��-���Ġ�z(h��e�00Ǵ�i�o!ҧ��0r*��a��)|��T^ץv�Q
Uһ���~%m�=P1�#���f�6J��u������3K�Q���E˕�?L�*�v�V��0����QȻ�|="�h�ɒ9�X�6��i!���=,���e���z/j��@�S���Tw?��e���Pz��E�tn$����4�tѳ����
.��FeG]m1Ѡ���}|d���Q`�K�s��~[%0$�����m0���2�,�;�5����3m�|��� �^����`)�|��c|mN��Y6Dؼ���{e�x�ݓ&��Ⱥ�W��w���ե�]�]5K��gS�,ka|���	�_�/�;����3,��>
�%X��&����D�:�@֍Fl2.�@JS;¥"��Y�B2g�b��	ك��KQ�����% z��{�P�����W��o��]����ʟ�g�Z�h	��F�<r,G��Rt;'�b�a'(�D��N��T#�O�[�%����K�������N��ސרv&�y��#��U)~H�Rڹ��'�u�{��,r;;5mLB�b��f�j��aǏѭ?�	��5W�A:�9 ��tȟg�,RE��E�!�������P%�7�I�B�NVJ���&����k�;��+O��P�c	�8��B�[+�#wf���������A��O�Д�fl#��/�k5c��u�&YsU4���j1
Q�k�a���5?�(V]Qz���I��{��Ft�ul�s��B���g��H�^2Z��\���l�yz�*���!�4�r綉�#Jz�j��V{� K��-qiX�r:Vr��"$�I?��!����k;[cM0�Ѫ`�z캦<����F*��Tf<�"5��K�ls<�z�$c��rUU&����n�c{g��*$�h}�x�jo������]O��(�_�	�x���nS[��9
�b�	x��
Qf�B�xkMsni��(��	���ˮ�b��3����~�?���<M��Y˴y�?�~{G�Ӎby��59�t�Ս��>���0�	m|FtiUd��9��Fs[�@Yg���T!Z|�͋ �7<f�Tu�eƸFӍ<Y}��f�����9��A�Y���m���n�t�)������l�?�X?�Tv?��2p�k��kl5MPP���,��n�@qLxiBI@{�����lU[��.=�����xL^z�}�NIK�Ó�b`���Xv���o
��,���ge������d�ָ���B��%+����n�'��Ǎ
�o�w�p.J/��cYQ������Mo��ŕ�`�џV��[ޣ�[�q&ǄQ	flfFwq�6Zg�eN�?�&�J�f��t���z��:�a{t6áx8H���8\�� Ϣ����O13ǜx������fK�u���|����0�Y��yp�����W�hΰ�A{���2�`8DA.���z�ԝYy\����^��)E��x��N�J�/I�ĭ��{�|��F����(,�	� �/�0[^��� �htphpxx�Wk�����"�@���D�H�{��`/%�)1�#¸-��w)�-�8گr��[���++�w�� �����kd���<�D],�m��,�q�k�s�\���B�a^�"������v͘�{�W�Hׁ�;��b���!�Y ڦ�Ӄ'�J}�ǆ�|,f�c��b�w�>��<3��;��;}�X���D9������.�wz�z�C�4���H'�OA��"v����iC�¡ ��fx�OI� 8��qP�W�S��u���������"�-Зk+D�S����S�Z�Wi��6Y?��ډ��c�_�5�.�q'��zfC_�l��8�������k�uI�8L�jh�.S����.TtO%��@�{�Y��`�ZL�	 F��1|��wn5��Y\gxP��\���`҃d|l0Ak�����=:f
؅�����i���SD���B��a+�x���_@6=*b4a�8��׏�m(�J$��Ւ�_��D�e��>�6�����<�T��o�d�&8sU@Bm�Uk���~���z3+@����\�FuR�o��<��*�����0Q�"zJS&��\��f���1Y�*k\&ڲ{�����h�ӷ/�A�zE��a��Nݔ���8F�\�H�A�7jT.�iֶ���rBm��}*�*�q\Q�dK�,Ǿ8/���<��ܙQ<�(���c�X\�d��ŭ�Z���	�R�D�N���N	p�<*1�pH ��+C��ke�ӷ�1t���Ǐ�tI�w�ZOP�!%#[�C�����	`%���77�6�X���g�v��D=�����6����މ�z���f�xp�j�:~�G���k���	ƪ�|�H���Rt-���W�'��P/I�5�5n7� �+�\�0�!��C�t��
�6��}oM�Q�K0>h�ݗeFx�(`؄K�ߊ�̺��_�5�M��&J�)�s �o*�Jii�?��#$]�K;�n�<*O�IУ�R4�Ll�Q�dI����&�a�X��b�c��k�IU��?1ћ,��[,"���n���,�y�9�9��R��O���߭:%�%�U�FE����hX�*��\���f?��Z���jk��D�~.�I(H������XJ��v\@�(Y�sG��I:\/�Amx	1>27><��M�(�ݴ���8E}��K��O-򰓛ד1�1����%�Q��M��OD\�ִ[Z�#)V�X!�5�Ƈ}P4��D�UHL�f3Xp�Ҥ���|�aኇ�F�A���RM��t�oaJZ��Vj�2��������#J�wb!c1/�I��Tl�<Ng���'ߌ)��
.�Z���7���頠5׫?��J��V��q�}	!��j��H�0�>­=��W�W����o��;r��Qs�H��p�G�nﲪ�0�!�DI1w��e�D���;��?�z���|N��n��Q-�_(�R���������d���L�I1�����v��Ou��8�d����jh(`c�t����� ��%t1ߖl�l��j!�	hU�|4�����xj�(*vI�`�u��%.�c7������DMf��+G�Y���a_�L�� �'@�� l~�b���7B�G���ne-�6J�b�]
��������J�x���\]0ih,'�6�����,�[��]~rĈLdv��Z�`v�;�iFO��&�_�N�����҃�̎��g@����"�(݇��QQ@
EW9�~5jBXZ�Q��y[�T��*�AU�|t����}gސ�c�Zf�@�3����:�B`�����p 	k�r��I	����}���O��}����Wy_�i�ҧ���4��=Y�Fe&�z�)z�#GC���a\U�ٮ��8���I�Mҷd���Mxf�p�H�R��~#���?c���e��?�����M�L�!�����P����jof���LHݿ�4t������ޮ0)��hlV�F�����߃���he����6aPt�Z��,9��O�҂9Lh�@�ve+����I(�!�7�ߕ�iMt#�y�i�J��Y(n��[��H��֋���@&:j�+6��()�N>2�3��7�r�W��Ym�5qwÇ���9������X��M�Q?��F֤	��H�"��i�_:���+�D���GMaD�5D����:Bs�}6���I3j�/A�XB��?���ߧc��;�O�$
��̖�7=��-����Q���")�����Nk_����!
�a�0V�,y��)�H�-渖Қ�� ��8^8-�5}D�<��`��Fc,����G(�:	�&�3APtBگ�;��4J@)~�	V�x���*$�d�R�͂Nf0k�'����� ���9Nf�F��Lz���Uzy��=f񦩚�,Cb��n4�2�մ@��G����{rq_2�|���9�1/��p�!.�����%e��Q���)���C�: ������H��Ԇ�ď唉B�	0(x�ѿ���`�hyeq2�A'�w�5Tl�yK��sRc\G|?(^@��J�?���ݦV�Sӱ�w���q�oU����j���\���`]���Ry���DC�,~�iZ�\��
^�Ϗ�C7���g>��a�x;��L�d69j�o1��T.���1M���hw�<;�ywL���c9t�ڔ��ӌ��A�_��N4����ޞ����Qo:$q4Y�$|C$��6��� ���;.�oEx�(p�H����r:���o����t%�0)����5J�AԠ��LYZ�ӂ����z���������smw/
16{K�
��9��io�/�6��y!��@g�,_^D�%_y� ��{����՟��������qՔ���ɾ<Hk�h��|+�q32bk�}Bq��U^�p�]��f�a��d�%����]6���ٮ�Ƒ�,�6s�޷�7k��8/.�J��y��|���E`���<�	����lK�^>�*j�$h���u�+�Y>�eQ����V�ã�ռ��Y��O�)��g��4v�7@�/�	9�r��X/�����P+��~E���ݓx��f�=�%�9�ŧ�Ys�wr����Ld��Ǔ]m�+_�ۙk/:�g�S̱)�ڿ�2	����`�[�h:؜�ng{e-�����Q��E����û���I��{r}��	O����،�R��h�;��f�uůٰ.	���{�n��	|��e�6��E/�}Z�Q�3F&A�(#�Q�$�6� '���΂�����Z�K�d���9����^�[���_����ۈ[ͱ��0z�dҒ���)��e�t��k$Z���Dmbl�9�r�0?2�d������l�<_?n�;�A�VN�/�cN�����{��� ~�޵w�z�'9Qe�l��fV&2����:=�m�ۓ{Ў7�i�\�P�]D-ek��UBԏ[y�����G�'&���	�,�*o���y���+���ko��s	6��ݤ��b��b��~_vJZ�҈�@��+Ui��h���d���_�X8�P����#�$n)^c�v�"SY��p�1����.$���vF*�v�{������|���	�53�������W�֐����o���̛�i���al��������[��ꏼ�?�Td��n�_�[��Ùӡ�م$҅U��݂JQ$���C�P��i}㩌��[Nr_��4	
[�7K�ɨ�������S"1YA)���W�uAe�nF�τ�ms蔔��lK��Z�`++O�D`5��&ev��?�o�dət]T�+
$�.~?���:��d;;R^D�c☸�goVDO��x� �����*�f%ֻ�d�Bϥ=�zA[�̰�C��N���O��ٹ|R0�.2���<�w���L������FUH/�xe��W��be�2��OD���yO��
�]���l/hy[dM��Vx�z1Kn��V��n��-?�3d���ц���b@�X n�h3���Щ*?���)�'4���Ν���4Tl����E�ddO- C&J)'�~Sn�B�}��6m�#>�n�B���Y������Rm��������C�n1^@A���f+Td���X�ZZ�!I2lZ1�CV]��S҆ŭ��5T�n?4�3*�>��^b^�W�7S���1�� Ũ4ߥ��	�!6�����ez�K���g�,��,Uw8��ܮ��qMm�6M��/���h4��@.����Bd1�J�re*�:��rz��mF뵧�Q�����`�Z�&��2���ggq�R�
I�L��+���T�~�$�I�,�iJ�F��������җ�G"Ża�T��L�xY��yNP�����
��O�%׬B9b�m��RtdF�(}��r�U�{Ւ��٣�v	�ok�*��4�|�>�_���k�:�<֭�C�11���l�Ơ�_����� Q�t#hÉ��K�R4P�#�Y[�,.!QVU��������I����l�(%��]��m.���?�F3�n(�D~,�?e4�����d_t�@ֺ�-�v��t,��ݙ�9����,���Dgj��'�^f}N��P{�7�ء1fb�;�p�3�bڸeE��]w���2ml��עY��&��f��/�JC�'�c-����l�g"ݼ[Nv`�C)�_���|�`*�_S���O\�������&��J N63 �V(�Tݖ5|]AǏ(Z�t@��}��H�k|���pCA�+e�MH�bC���O[˄��b��]��>�%z����Y*�I���I$	ب-	p�'�,�'f�'E��{WǨ]fx��ֶV��"�q5��L���
�d�h}�&'�-�M�7_klڪ�1��D#�o�/c��XcMZ����H3��5|�e�PJ2��8���W���3��I�i�@J}f�5�������&UǤ/�ꙵ�0�F�*�WB ���'$���j*�G@̤,��;F���<�\��E3@�`�ՠK����v���E�W�`j�Iw�b�&I��q9M�f)(1����0G;�!��K���џu�=)IG�<����%��Bȕ�CЭ �X���~�/3�������.wzV�>�v�LW�]���t���X�,Q�L���0�D^R�v:cк��'��톮��Z���\Y�I�EeL���Auc���UQ�˚�`��K��h4.���Q>�;���A��ZN��ć�e��yk�&�%�$��g�x�=zxg��-��/.���r�Z���N[~s���l��a�.�u��_�l�O�%S=IDm�Qu�H1���(o�͹�n�p�T���@���� y��L�[�p4�̳������������O3�!��}?��ι�G�*m�QAu�88N|+�/Y����)� �[}�1+�ً��O1��T\���jN�pȏ��L#���h��pŧ�1�}H�Y���Q]�r��"}���8�T�eF�����$e�����Ԝ+d;v��j�I�+a�Hj�]f2(�����3`��iFt`�J��#�ܬ��vς�������K"�s����K����6<2��
�?�H�$�t�iQ��
a`bgU�㟗�n6y7�"A���-Q2Î�;,����|}��_( Z1 {b�Z���VP�%Gè��|eJM���X U�a&C�݃o¢�"�ҶC���Ġ=-��tf�H����b ����A�~�51H�����������m�~6^#��rnl��!)�J'��1Ԩڽ��2t��b�darśqAnS��i��>�Js3����Z.I���gWD���q���12��?d�FI`f�tz0�s�;�Ac�\w���a�ݧ��4�w9��R�	G�-���L]9��^�#p�a���q:�ic���=q������	j�V4��.��:I�o���X �����0T��
eݨ���:����W�Y��Д2G������U�{Vꏓ���7eݗ�X�:R��NRФ&K��n��RF��Ύ�֕:��5��;�:"��E<�TGgy�7N��kӯb��^�4_F%}�Ԉ�����y�@#%f��1��J�Ԫ X~�����Ò�>}]IY�Y�����=��}�4�Èt�P���t*��2"be�b;��*]t�OT*Ʌx�֧gY����'���=-ݾ����Ne^�>Zf���=�<>�բ0K�ؗ�S���v�vA����c&�ίrٶ�OŽ5���vI��ia ���_p c^�Z���������u��8xȅ�;�qT��SW�]�j��yh��f�0p�E��f�c���@AV�����l{D��4g ]i橴Zv�[��ӝA"��,.L���VՒ�#T�� Ơ�?���*<�8Qi�_��/�X_z/;�H{.q@=�	)M�i��7j%��<=�k}UO���N�{�p&$��������U$a2p�pG�3LPn��.���0���e�k���ȑ�$2BZ��T0��2�_�����V�TU�9~��;W���� Ĩ7��y}�5��>Dǯ��P�5�P-����>CL���w򃋲Y6I����!*�L��r}�q
C\��VT�]�ݶ��ϝM�Q95.�=}7�͔���~J�2��%=5��/�����J����D���zҳ�"{`{��.��6SD�!�UI��߉�~��3�J��"͌��@�K���)��^�v�Q��	4��4X��T�T��X_<��rb�2ujK�֢� ��������P ����a�oq��;�KP���D�6i��h�~����X|���sڬݖV��f�i��F�ɭs\��Q3�aş����B��*a&^?�|�Yv[��B��>�p����ٵZ��n�.l5�e�-}6w�8IkH%���w��������am�)z��~K#6� �y��2�CgGd&K���r�U�>Ǐ�[���
�I�ʢ|��VE 9���K�����H�z�i��$� ���aA��L�0�J��T|��Q�b4Pk4mnz��Ė4���	 9��Y4'�=n���tw켎��$ccA�O*=�R�&85��i T��&TaJJ'��N
(aD%�	A9Y!�c��0�/%G%25C��R��W��8sC롁�#���X�\����w�߫rjS��hh
�����Go���7� �J�Z�q�ꋅ{YPL9Z�r��e/�3F���?������*Ɉ6n����A�^�*	+b%o
�p'���x%>�(z���D���w��+��+:�*F#i�3�J��b
Kı>,����+r`�T�ʿ�#@�N���4 �9��	䦀]�c����{	��(4
��6%�Nn%�c����P �!��i���~D�Gޮ�Z�ōL"���	ʿ�����	:0F��xr	q1a�v9��6Yi����ɥ�a>̕uR}m��ͲwH5�ּyR^���a��ф�hmH��77G�_���U�\�������]m[�NX�cV
��O��OA�tx�C��Ƴu��ᨻ[�_��|�H쯠(;�w�!�g%P�R����@��,��Z����s򾣙���^U�|� �c�e�/��s��W���:�֟�3?�AD7���F�]/����sd�%��ǹ���ɢ/E /���vlr"it9�����Vh�I���[���w�֐��!�Kό�6��ۀ��I��S���L����
7��+�ɿ�Y[�q.�_"�_�*���:�:X�f���>$cu�:��֩�����f���x�喯g�)~��/dS{���uWSUD^�����W�}�n�K���q���4�&c��!���߯K6LMBZ����[��w6�&l׶8Xn6�P5_�,�2��P��MX�߽3A	��&�?���q����-�O��9��'���i�6i��ۺ��%�k|�X�A���.M,�e	�����W�=H!Z�}��1=�I�j>�*����zP��^�WN���v���ei�b��5�5�����PI�u����=w'�u)V���D�0�ŬދF����OԹ����d�j��jI^�&���jv�Ni���4�G2b$�xr*O���~?Ȣ�`~Ye�`��bm�g:�q��P��:ۏ]�����6K��L�,:9���Q�aB� .���/g�����0�B�h1|�ʵ�Ղ���-�d��sl����kc�oki����9�!��5�X�� 8r������a�x����vGa�ㇲ�������[!�,�^kٳ����ih���LMa�n�F����L��Iy
6��j).� \O�	��wH,{CG��*:$bq�L��S�]��Bb �a��K�b;��
]b�"�a��_�a#-�Jvc���Q+���gsem�\p2��y���U3U�F-�i���.�Wr��ҡ�:`����r�_�Kb�a47	M�	�wř�r��W�Ctp�e	��t�����@'/��7Ɣ����=�V*�%'t;�����K�/�魕]��;Q1�w�jm=��	���U��9|���Y�Ʈ8�{���"Dd(v��A���t �V�u]�j��O�2迾Y��3=H@���' ��Y�a��L�U<gc��̑Ho��g0��"��=0�Uo�����&-��?��� ��X�8A�4�Px�Z8�%v.1��̍�ml��6������R*�?�[q\�xĕ��N|k�$3�zbtV977wbjJ!n��B����͝^��jAAN�}�;�q�{F|��x8o���p����4]~b����.�V�������N�z�cc�nR�H�](�]z����=�M��` {/7t���>$�$�����F����q�log����9-�BL] ���qf���b�P�����%�����s�0 ,�f�g$�[�i��A1u�%\���݊��h:�PR
2ƀ4�t�8���âM���39Zrd�0�Z�5 �B�L�?і��o&���L��g�n;t]�lY��a�:�L�^�@`ԙ�ͭ 6f�_ʅ����,�~�����O؉#����f��Ԑ���V�QC���܍[�=1�	)i����2Y5����ʔKn�/�t��V�Hk�Pw6Ar/�z+�aĞ\ � �a�E���: �ݵ��!~��A��1��ԟ�@N�Y�r0�^����,�t�T:���o�a{�hxX���A�(�vo�	�bWW� ?�ݪ����ɮ��Z�T��������ϲ�0+�,(B�b|��+OU�_��dmq��ɔ��rF��j�����w���$�u�T�}:�;7�F3\׀cV�=f	�r���^f�>�-����ڛ޿R7k~8����"aH)��ՔL�d���5�_}��I����\�2`�ըhߛ�*lQ����cb������i�gk�"	L�����ʏB%eͶ������GD��,�`h�E����ݑ���Ą����L�q�$,���wq�
�ϊ�fy�����j��𕶙ƸBQ/��|�a����E䠮J�
�cG��" ��H��k��6�J� �������j&�F�6��V��̜�vA�r�Slh�	��բ�7Hxh��Աyk�s���S<��� 2�X/!�+�F�ޒ�ùq�qw�2xA���	��^���C�����^P�+�0U�1dng>��s+�V�~�z_�H����j<�ph,���=
�ط'���7|{�`k���a�U�}@@7��8�Vr
+����	s�����L`�j�(��!K�:K���զ�G�"&����w��!�$e�CH1$	N�%�$�r�'�V~��ٿ����@9C�_�5�;}eS�s�7�s?>�v,p��)�>��T�A�6�_���ɶ�X������	�����o)�L����'X /�|�6��j�եn���SM@s.m/�6�=(l��&�_���Ӟ�u�r��W}`��i�"��UA��2�Wt���aX�D��T�T�O������d}rg���~D��}��pV��$X��s�T� �>UAJf�XEձ��ܰ���$�h"ɦL�+6<n���x�KNr��ח\_���(� ]�P54�oǇ���~�ޏ�4Lt�"&%|R���՗9�cy��^�>T;D L�hH|"?L�&F!����A�۲�O�	��uk7�[�R#,�C�_@�v�&F��R�7�5)I	sĆ�S_U?ي1:�����%@�E�\a�iWo�rg��X��?�>د��9�"w���XM��u�1X��%Ǚ���9�U��*�~�z�Q�6��!�$�r��A�z`�ڀ�����V�$u��X$�n>��-v%�~��3A㗕�����%Z���k)�;�S<#�p�a�Ϊ���"?d(*ᣴE���z�^-܌��M�����Ɏ�.) ��I�bYit\)�JP_c'1�o�k�	'�����VNY5E"*��RJ��TKz�l��=�糡.�a���I,�P[�sg%>{j�r�gcL�R��ĕ#�����t�w$e��\Jl�.��o Qu#iӺ��{�hH��F��6TՑ=�醋8�z{��\X���Ԉ�J�c��;JU���+��V`\k�#��͋Y���Ė~�,T�r����=p�Q=]�Pz�]W�ns��'u���ڟ�)>p:;l�ԕ�X��"֥�K�N7a���I����:�鴛{��Q���7�䵮��[��C�
���ت2��t䓩�ӟ� L��~=:��]��[�����H����eN��}�x���YXM�\�*�8�W�*�s� Z������ΈMՔi�L*�Xl�'
_k��An���i�Hkϫ�_�X�iܨͻ�Ữ�,}��������5o��y�K\xk�`�e�kХ��_�ǟ��e"�9bV���uJn"J�U)wq�5[�es@\�YY<W{
aU\�=V�������<�nUw���HG��
8E�	�ڟD��b�NF
����ݶO��eɟJ���i(��ȴ�4�]`�-���/K��ʾ-��Vax�e���WO�`������� ǄͰ��sa{;�3-*d�zI�+z����2����^*�t�_:��{�]����2�Le���bbK�v���x�OW�t �3r�OZ����� �Ǧ�.�o_b�t]?Bխ'!�+�<��U�
\�:l��6�9�݄d�br��'M�8����g}*RD=585�� ���]�ۨ9��P ] ���~��:�P,h��=D�c�;������cs��s�����Zm�gMd6�r����ؐeLݻ� aτ!�$�)C,��$y?~��wt,��QI�M��s[���5[�t��:^'� E�/��,������Wl˃?i�����G����@��C��st
��w���/��cwql��X��unK-�*ܐ�ژ�� �ѥ�r=}�Y�zn:p�L�W?]ʃ��Y�Q��_����(-����~��SP�$���dԌ�����e{3�s	�3��~�2x���K����7VQܿTo�$�1��N�G-#TPM�������F,���d�4��\m)�b���Q��U~�^?�G}l��ؗ��S@����K��� Ƿ�����T.=A�����i�UmO�R��� ��X�\�]Nӈ���z����~��Q����sD�g��3�����y�>��l<+���r����a+�l��&��/n�mXoS�e�2��;|F�p�Z��E������+�Um7J�*��fh�'�#�p����E=]��开�d(�ej����Xu�v�ݩ��x������C�V���D�A�C����]u��BR��^
������밾�oM�?#&��<u�g�q��N,\[wx~�vSY̱�w�,�R_�;k���7ŲT؎/�B��c�"b_R�@:Oq4��w6�!^��� ���qr�k%n�J43��Ӓ�P����r�\P<�3� U��Ⱥ֦��'�<�3��p�.��t�rһ�?4�	C6/h���y�x���$}��-�u�{Z�eﭤ���ӽ�_Ԑ�/Q��}�7��������E����Z���v���������v$�s:j}��#�k*N�4�2nbr�v��X[�ߩ����E�G�E�'$�L����8�Qc$Q� �֫\k����u�)()'=W/���m��Zzl���GՇ��`6�dU��r�NU�V菭��.mn..��
'�������~�S�q�z>gT�.l�Jd9?^�J������>T���ZFo��쯰�F�΁G?^���)+۵��2`PJ͐8~�9U����gT�#�3kj����|J����K�k�<q���v�<j�rv{T>�o�q��}3<����P:'��:����Uu i�sy4�c�,�� �7��^���̅h8 �fU���伷$V0x	u�hf���O)`�Ѳ>bA��̣�������$tjg��Ɓݩ�+�MU�J���D��ї�(�ދBs�r<��ϵo�ָ9.rf���7��( A���������7��L�'\�5�Q���ֺx,���-X�	���{������/��\��m�_�~q<@����-��Ȩ�B��`J�*��)�<����;^x|M x����5�=����	�}�?��^�v\�Ԣ;�޼_]tB$����(�}���j��x����L/�>��Ѕ�"Z[)�(f�2��u��K�TL����-�|���Wg(>���s8W"��۝Q֒�;OH�CF�U�~t�7�`ۊ�����y��+R�U�@��d�Iٻ`V�2C����ڊE� �\��q�=�Z<>s��}Ò�2.I��&:36jZ��o8��wW�qV��7t�J`	�֮��gv�2"a2���,^��8*_f)c��!��S}�sZ:�}�t�Ѭ�I�ےi� #��n+�,��`@hي\	"�0kS-F�L���0�G-2Za�2�S��6-7���U�zP��#sYr����?]��#7���c�m������?F�/̹t�*�A^i���
;L�>���wi��={�g"����3����UN�J�������o<V���S�p؎(��c��TAo�Q"�Oq��d�~�"��O7ș���ŕb���=��j��USP� ������=�|PQEu�Ӧ�nܦ_����1�@C>���#�d-�y�^M�@B�ܺ���I|Ͷ����Z��)l�Y�m��LXr���<xL�v(�Z��`%�����QQ�_�(ݠtw3��� H�
Hw��tw� 0H��CwHww���?��Y�f�{�S{���sY��Gaf��j�cZ�I)*���ki�g���(ɳ��s���!o���LF&%=S��D�/�?<Z�T̓��5���x=�/M�}ݼ`b�ڼI�j?�l�v=��{2(�ײ�w�Cv0��
S�8��l"^a�
�J�"�}oSf�c�Q �����*�QC�V���������T<2�v0)���2�$`i*Ƹ���H�r����'�I�"�!{I�)�����9�V�uJ��������2�x��\~�:�Y��*�WbD(F�a��F??��&J���9O��1^��6Y��U"��N$�����}�8��]p8�-�b�Z,i��W���f�x��,R��2�G�v��
#����c!��б�q��½�Hߩd0�"��k�6K�â̩i�?~���(��o,��}*2\\\��Z]�B��}m��?� �Q�#@�<3sbvV�����k��1U�g����nq����t5��u�b�Ƙ۶$6W��G򖂺x�K�k��09��E�'�p�wo�b#��8lB�I���@�~��M�ް���u�͐?u��x��Ԕb�]R�>�+�Xօ�P(�7����:Jj?$%_ƩWR�y��u�&,z�����@�dm��\΃?H��ͳ݃�D?�nv���]Q�ZO}�����L�ˤJ�jAl�Ψ%,�Ө�[)��Ɣό^b��☩s�nm8 <j�+:�p�t�^���d��8�ON��`��>B�/�ux�	�$V�m���~b�]�]�1�&VD�|"^EC(�+ TE&���K�������sLv���<��p�47����=�4k�����+ 
�l��@��*����N�o��U����)������!VFSI'��oD6�f�(��LA��_�Y-傠22���P�exG\��+��"����Tz�G���ܤ+"�֬>3��Z/�R�//��!�2���ڨE���R�$�;4��. 6"�Կ7N��_�b �C�'A�Os��DC_��Iߋ��!
�_�p����hoe�x]�nx�$��0��M���V��Q����K��T�3D�
^yӥ3�3�F����`����T�
�X{��*��|�L&�>����%�^�_�{�jbWp���?�� �F3��0��k�)X7RC1���<K�*��9��>�����2�S0	�ٲ� 	������FqN9�y3��� 
'&+�m!��clc&����ݮ����:[g�m��lI���,�I�� (�WB�?��rF�Ⴠ���J�itj���?�I6���(��R�M)^������Q��33Iu�0.�Oe:},h���&@o��80�Q�5�\e+�`::��%B}���*jP�~�1UP��o�N�㡆�6�F,	�	�=ݡ�z?��T�Z!a�Їj�ڣ��ur��!qB	�d,��}5�c�U�Ē�9�\4�)HC�A:�	)Ꚃ��2X�X�/��q7ǖ��^O���?�o���li��b���t;�/zu��cL��%s�"�����&`(�ޚv1�I�Ol`P��r<�x;Z3-�3!��,	H�q�����5c66>#&^fr3JP8��0��=���(��6���|U/�Ȭ��F�s��C�*䎛(`G2���|�`-D�L}9��	����������-&v��S�p���F1S� ���D7��,h�I�+���U({u�8�nBN�8c�.NP�"�/5%��U����f�\L�DC+�%Sӌ/�k�}(��Am�[�T��ɘ ��I��N�p��BC)�d��a���V��+n
��^-�A��ơO�O_����{���Ag�,��������hn��c�ij�f�]�!P�ߎ���ĬjhGFV����6ʁ �i�[�A��Dy��}��3"���M' ����y�s�.��l���(�ye��oK�C�8HX��׋�|""��U��ϳ���C
.�1�K��HR�����\qn���f�"ڙ}�H����l��.�$n�G��5+UT�� tl��v�7q@���JW [Z�wB���ݑG���τ����^)�n�A\u�P��F'4 a���Y>$�_��B�{8u�wZ� �o�^�B��B����
�Kj(���=6����}%c�_�lq�ia�����V�:�d��(�	
��
R�珟t��!�����8�RA,�b��^kh��E��+��j)�b��:]�A��Ȇj�QϤa�}�3�gby���7�ߥ]3�Rت�C���<�,{�ow�]�><��%w7l��7�N�u#����o0m/���\�ӳ��/Z닢�FvT��a�2+l��^
���O�/�����|`���ex����/�cyl?�:�vSR�n �طw����Н@3��\�8����>��Y��l������q��Wk�VSJ��}�NBR���N����+q����
�-��3�H��D����o�~~�u� ��B) N���!Ji�X��@n�l��!c]��<.Ka�	P�F�:
��8z�6u�(���/}�BB��sfzZ�L�*7����s|MOUr��̻�`�c��3N8�J;��3��׼m��Ԏbz�����
��t�Y�8����sE]������ʄkF}���O��W�g}ˣ�r;E�7��U���M[Y�%�eE��57{�.�(�����P=]u���s=�\���W�I��k���X�ܫ��-���"j�ͯ< ��~�3Z\X���	x�*[�>��xl��M�ugSZDҋY������:��+`�y����1ϣǬ�93�<G��I@�����������7S�~���Շ�9J�2��~ּj'=�����.8��k�['���@7��gl��s?��(y��߀��>l'���L�E[e�4�A|�x���)m��Uږy۽���ά�8���59[m���G���ZU�_���,�D��6���/2B��ˎ����dM[K��%%
�N�8�:��񺺦�u6��s��U��ߓ!��s��«�#z�3S�-�B�ġ�Z:W\��R�e�b�.�f�s�r�1��s��I���?�Td �9*�������6��C��v��{�y5�?[;ɞ�|�{{7ge�Y�G�)İ��b��s���J����Wf�����.٢�	h��JP��C�4�3���Q|��q�SO:DT�)�ႭoEӘ����5:_1�X�Nb��ճ����s؞�4Q���~I�9��h8�K�FcM�/+Púnd������x-Nu��Eugw��ҽŸ��Qgc����fu΂�_�m���`ae�Y5�5�)	Lx0���~&����E�e���-�
="���+r��a|)F��C��/���Ej+kg�GKe�`R��u�ۋ*J��p��/֢��"��}��Ζ��āGٺ�Dd
�hv��^��w�v���K?)D��C@�d�v(���~��c���PU*P*��d�l���q�����$��&�[�!��+� un#�k?�r����B�{%2V�)����e~wHt�}���s�AQf�ˡ�4��5���1��U*�ơ��ma����Vi�Q���r0��n��I�Z���\z<�­8St��G>X��|�'%"��p�T54h���5��0�D@�J���+�}�If*=;B�h2�a1��7J��Y���do4�����������l;������/���J�vL޾B�8k̈����P�4���u���&p��⑅�V�8t�3�UZ�@-��>�;$�_|�b�x��s���0�T�����Q�8\��Fy:�U(��l��Tw�a�`Ҡ��}X��,j	u��x����'l?-U���׏��/���Ԏ��0�D� ZF�F��B	�0�s�L��/3�y0�]�s4�<��ъ��+ƋƹBIS�Yሸ�*n�7�<�׬�,;����9g��,���`��o��9�2j�'�%�C�)�>_&�+{Wluh�e{�+}�p@�Q�����-?X��"�Q9-��nO��h��U���={$?��o}e;��n��6��~�<��˙<��#JoX��`J�������Ӱ�o��q���,
!�m����+���D����gNS]7��}�Zrb*E2��q�v���T��5{��9n��Ԣ�a����a�C74����5)�W����}�<<a�8붇-��O-;���?��1����9Iڋ!���N�n��4����%��?��87W�����跙0��}��`w�m���ؑ���g�� }��.���Yn3EtF�^˻��gL�<kԬ�z�����#�+(��,	�����j�#Љ� �ha(E�'�BP.)���>�da�H�?�oQ%��n~��ru��N��C8Q�ro�^5�~�mi���E%Ci��#;��e�0E^���M�D��^� ��׊���
O��*�,����WRX[φ=���lK��$�|�,&�>F׫|�o7�&�riU����rĭ�t�0�p��������#�����P?X��r����c#�T��o�DA�1�n�����Ӧ���B�C!��:���K.�!h_�Ѿ�:>T�>*g�A�>�|�$�K��'��B��=�C���ss��N����V�Bf��:��']�҂Fy�w��Bv&u���͗��E��mν��:�"Ӵ���]�.{���oZ.����
��
�=��$C�.���G���1w�S
���ˌl�S��!e�t�?�_8����WX����D|a�-�}�* �0r���u[�6y�:U����Э_İ;�G��m.�	
�YV��DQ�꿹{xޡ����l���Ʒ� �qA{d n��2.�!	_�~݈��+��|^��z?F�i������<s���\���%|����h��p�����]C�?�6!���)��2�w�w�1M�u�v{_��fZ8��<�w?�,]��WN��i��}�>N�ܦl ���&��dR��!Y7�m3������L���xį����K��xVm�+��;]���¡���İ�8۰�m�Q��w�C��(�J����]Z�/��H!ުu;6w�	�LQ1����\p�`���!2�?����{�?8��2�۞���wNz�OAW3P!�Մ8tb���p�ԓg�Lg�U<2nc��8n/��fP{xz���JCe
1wF岡#XޕJ��8>3+� �W-r��@+�3�^���n�i�<+Y��QQ+����a�f�q�A���%���VNu�z���,_C����5R��I'�|ʇ��W&7���r[J��S�z,�_8��.'{˜����k�p_4����@n>�wХ*����SXյ�K�*�-Fy����8��H���c�B_H?N��Z�l����&R؏�R@:Wp�^Wn�2���<[�P�r�[����յl�gYYx����ʂDV�R���ͱȵ~d�}ETp��=���R�NR"�eH�b�V���c�۶&�**1�s:Uzsy4_�Gx��F2[�.�EB6��ӵ9��I��	j8#-z
���=.K�v����������t�؜�����b�W��1�}d�~�1v~��.Y&bӅ�6:�r\<�e�.\�m�	&m��^>���ʶ��i݋E~���KGÊH�i�@�H��\�Bq�1�*�Ͽ��]i*�@@���.�ue�w-��v���B~bg�5��C|�v�0�X��H2�RC��C���ipt�z���s5�l�����aU]h��H�Q��Z�a�~��n�ӨhW�٦���S�����B����F��`��t�^��}���pp\d��h���Z�{�@�U��GvvV��6��=GNx8g[n%�AS�s&�V4�%�=�s˚�X���!D	�h����F�ey��g�sd�^#5�H7������EA�Đ�c����*U��	���ٵ5Oc�2��;����p�+��PD��� ��HLY�^� ����iK¯[xlʕ�kA/=2�l���l�dĹ��
��|+�i�m�5kGّ�%�V�A�͝�_ڟ��_��)��A3֍-Z��m�9��K3�x��$�����{`�9�r[�2p< �%��!��~��������7ߥH�����}붿�"�C�~����Wd�����׳U�|^D����6���Ϯۢ����-?�w�]��D6#�kvL�r�^���G*Z�QN���K�����!�!�h<E��X��#���a�î�'�����>��u���:�˳�%��o��Ө�ߎq�d"dR��K����%���ﮘ�?`�]檋4�3�}o� �-P��z����&q=�>��J��I�3$�A|�Y=
����[�����
�.��	meЀ=��Y���[hˑ�?~J�Xn���t���z��{3��S�Z���a��z�)��I�T�	ރB��p��፯��m@��� �L��2�C�b�O��=�|�|0z.$�:& ��6�f�} �y,�x��-/ָ�������e�6���d���C���5�;6���Ka�9��rGǺ6�b�����]�Y�/z/7~L]��y>��F��n߄�[��Ì�ϓ�ձ��3pO�
�bh�Z:�I-�/=2GF��3j�;�Y'�|O�"؆2J6^7'c�{Eώj��t�=���k�����!`��n�����JmsUj�>�1�Q�X���췹�5%|��W(C������[�ۮ擐p��F�0I��cP�@�=#��E�7��i��Cr��n<T� ?�
W��gZ.��jSb�O~Xd���A�ǬF��蕧{��L�E�Y��bW�\��m�7�;���$�'T2T��� �BJ�Z$�OV�`w<F)=�ִ���Q�s��z����=�1gڼ����c[~�4Ǉ%��QzK�P|K�d��\�:G�}ik���٧���n�x�FS��sȶ2
�2�ma�٦[a�x���������g��S��XZ9�3Fi�5^U������@�0�;YY0G�ռ ���r��e�������>�0����Z��,�Uu��uG���pa`��aD5��1��oV��?�օkUP�)r�.�����Ց&V��o�b��;O%�ᡫ�g��I�ws���xx�B�E]�@�K(&�S�t~1�����+$q^x����';i�E�X�c�����{g@ �#O�{�*z����ۻ�N�׀Ⱥ@�2��^2#U�]t�1�i�&�)q܄�cՙF��J�{��+����Z
��}��co�<�qh���z��'���v�������*nH��{��\/)����j��Z��fT5J=j�Zlڧ�~�ٲ�>���A�>+�*l.gWh-&�D���Llp��5���67�ځ�T���-(XL��2��7KnE��~��=�@��
{��q��b��(�A����s � �2��$��� {�A����{x�O1�#6"��i5���ܟ߅��3��^�#Pd%�T���fK:�{;!>�4�����i��
"Pja��Rlw��B�+,��������l�k��7���# ��A�e�Т�M�ShJ($Z�L{ʘ�L�6���~<O���&��o���}^� A���^�̝��@�	���l�E���Lž]K��_r�V�A�I��R���	�/:nW�[��nE5>�����`����
_���ƺ]K�'^����ֹ�%���s�Ā�j��=Q�h�N�-�����fu�$ʂak��'E���i[Y��{����70���T���3�J3/�����ԢL�I�o�6��i�wz����߳��wb ll���+̯[����VLS�c}���o�Y��c�����jj�<D�+_���F&|X=�G,�-C��2��t�aSp�%��*pe�$J�e�^�\��T�rXIq)7��{���m�WH�[o"R���(W}�2I�$X��. H�ۋLtrʶ�� �]��G�A�d���fs'%�p�uP4Ƕ��j��S�s�~�_��M�u.�}��l5"HÁ�E0�F��ŭ� ��u	Y����`\���\u�9	�1Χ��g����ގ~Z�D|������r01:g�{��X�s�y8�'t��"�!�H
8��m�~=��(��u	��HN������dQ�%�q.���_��z�t�����u��4.�:�M�l����_�y��x�M��9w,���,YE�uN��>���]����(�@��Zf�6[W�� ��v8��բo��k��T�����/5���T����7F�?n�j��p`����b��51���@�wu׻g�H�?�x���#~O���a���c����_�n����������2p���&�Dg���\9\֩�NƧ|�y0��/��gL�~��
`���+��uD�9��V|��R���`r	�M�@�J��<���=6W"�c��'��E�)Z��!KD�~�:���lsD-���_��cr����*�=���a�s\j<;��h>�~/��FDP�ZB}x/���p�=϶�훗��|�J�(BݶU2�V4ԇm�-fq�Q��#5��02H
<�����4��2ou�%ʀ[>,Lƕ96���τ��p��f�\�����`�I�JWXO���o8�7MFJ�}���9�����&N���lTZi�1+D�J�eG�f��!d�ƌL�hZ"-�ی�\�4O����֪�T�tT�Qn�㜈��~���U&=�jU��G�|��6�ל�`o����~�681F��r�c��/�]���&(��/W��»^�o�&	⃰ȇ��㩨��uip@?V�P�zS=)��V�"���d�^؞AǗ�v�U�赜�_�.��6?ڨ���)�1�{��"e���?��@A~=Q��"����=G�DG�"X��ڹ P�5�֚7>��}Ⱥ$" �֐e�����o�ׅ{6�����^���{}hΩ�6rL*&$1@����|
��#�C�K�
x~��*=�+z�uyb0�9����!��C�?qS�V�µ���%!���GeS�XpPtS��0#�^�0�q��N5��G��)d8����BI�͡7Ϭ�;�;�����i���?�|�%�3�M�k��e�}�������6��Z�:�1O�q����oFm����x>'�=��)��
A��-&S̹ M۪�n����Tb[ P����(���B[C���o��r��Xs��g�i��J�0�� �MM���Ϡ��,G*�y��<������I#�Ck��' h&�+��x�ɢ���
�s�FeB,��4zu�s�S��(�$杴����rl�����	�hM�/�d��N�D󵞐����,���=k53��Ǎ���g��0�(ӕ*���u�����v�5!Vk���w�>\�GN��p�sP�"���{���MQ���-��*q%�~�;��p�D+�lڨ�(Zw��/x����	:X*�*G��+���ӵpV��Jj��{G�de n���'��T��'2JO�r�ӫE���,=
%2cz�������U7]����2#0�����%�}���݈P�c֨t�)�w�cdt���ʶu������V��K�R��m�[F��dОDGA��B�a�s'
V��Bw������G[�)�����<x/�wi���+w�fZ�N���<���O*�5�z�Q��O?3ǿx=A	Șr������J�jb���f~�� '����_����$t�@���7{x\�ٳ�DH�,���D�ZBMu�V� �̹�����l9������*���~�Ւ��hx�ˮ���ch�Y�M�oe�w�+��s�cy�)k0�7}�!�?�����u�����z�E�R� ���J�wA9���xp�&��F>�����Y�lz��P�#<.._1��"��Y����}24���n��5�P_���		h7�
��0��9�88��Ev�A�������h����o[�h����[�W�ܫB��vǠ����1�):����k��$��}��9�Nn"1�dp�1���>w_Ʀ��6�4^��qm���@1.LSpw=h���9Q�|,Α? �s`����L�뫔\�K�ߘ�����d�63n�O��,���������T�;�E��edK�.1��lf��,zJ�f�ݣ��]�^�$�|w��pſC]m�lFl�(l����y,��|4��H�[4�B����z��L{i��E���nD010��o%��t�7&Gtk�$h�9ˑ�����f�#BJ���n�-[�������t�7Gv�'�L8���t�ڷg��4��/Z�0+S�C䩌h�����=>�!��^��!�r�˦O�9�'nᚭ`g�v�.37'�0h�]����LG[��(����`v@�a��p�)x;��b�?�����p�T,��?�>�����W�LQ��kM�����^K4p�Ͳ���1�*���X����=��*>�^@5 �B+��:��b�Ux?�IQO1���&�^�	K�up*�<�a�����h���r�)�7�1�����J��=���'H-�v��"�)F�$�;h�m�DC+*6���q@�ʷ}S��GD��ag/�K������(<3��ψ�=2�W�M��t&>��;Y,�^p����f/��¬�֮<	����{l5~���/9�.�(�W;+/r�BZ��!�J8>nX@�^br@����P���-4�>���D^�Ж�p-M��%�0I�?#m<(!Z`�#�%����jȧ�����	� u�L��UHɞ);�-�r<�C�:g������i��T�� ��2��W�H�&wCY�侵���������5a�I�8\�s�:���?|�M�I��g�*8<0)Q�"��� #:���sO�- ������؞�dg����v~~^�U�Z��}�U�,0��~}������n��D�7��_�a�����Ȇ��i$�|k����-�W���,�Q�Ұ)@�,������5^����Ѹ��8�0骔�6�]l�,qd�4q��=����Vg��C�q��~Zj�$�fIԪ��;�P�u�\�JbK�r E�g�.�@Z��ޔ�r����1��p�1c��\�ЎҮ�s�T��w����[ +	���mI>�5vI��片&���Q�e���E�"E�A��Z0�0��|�v?m���������|)�Rr�LM�./��u�M\-6_��B����5)9^�3D�&M"���V�˞�K��2��~:O�m���F��BZ�`h�F�s2z��O�������a���=.ӲxN.T��
�����r���;T'���6��:*޺b��w��s,�4�%K����
c������IC���A�RH! O����=�`�ޢ`�,1�ݵ��"�C^�	ݒY	���$!RFH�=��������%��&�['�
C�ئ�����* �Y���[<4px��¡"0��D���h�����y�r��U&�|�5.�����[�Z�~�0's�X�(�l���|��A"U����J�%'�K��F\�-6��*��W5���Rg����,��3���+�K�����!�ϑ޵?���n�6�D�TS����� F����#bm4�O�{~%����P��pA.@���p�}2X1 U|��׀�l�⹓�l�x���.��������A�#I�V�NCSI��Ļ�0n�/�^L"��;�1`7�+^!`R�|��4�_�5y]��.���/���>���8��*��������[����G��U�#T�{�.�fI�<iۧ���r��[gm�q�g����&�F��N�* @��.Y"[�j�/��J.i7q��5���$"��I��d΢:���DV��U���O��z�J�� �)��PI��8A�LQ�X�=�S�'��\���Y����6�_����aV��qI�F���Ɨ�Do7@e�2��l��Ё ^\���6�/�Ƙ?	^��Kq��`���t�����v�n�Ol]~ˎB��������ס�[���9��3�?%��V����Ԑw]���:��c��p~��KY�j�J�g�vtx��u�i�m	_�-n�+�z�m�.���6��rV���Ѩ��7m��B�8m�I�nX#8�R��T�PMw����9�b���p>���$��zܿ"�:�=tm�З⢢�����2�)�!�/����v�aSx'0��*��+>ѓ��p@1uV�)���-����"N���^�r/��W�n�2wO�Yy��}Ǽ�8oLR̮y��F-i�#�[�����u�.D�.g���~��C�����,�[�`�˟o�����ў���i�/���ߒ��שJi�w�pB�
�zѫ�<�~B`� .��Gj#ߏui�⦺��S�Qώ�B�k�hɻQD�OC��̂���>y��^�!xV�/��v�v�BS�������(�~��5���
'�i����T2s.O��m�E��fX�|��'��h`^b,��>%PesUU���#��p^�q,�(��v=���i4������`��!b���/��`�S���dt�x������]�������@�Pz�U]8C�L�wl���u����w/ĂZf!�u�E\P<,U����C������q1)0i"������ �AP����ni.nv�8u|2�L�Zu��uO_w�ǚ�z^(�5��ߖ�	+������>;�y���o�4�`G��l���G�2��8��LcI���D >�r�����P��.��ҹx�F��$�T1p$g����q�5x�����>n����2⠇�,��_bW��J�p
T�#�o�H��I/���ׁ�t��A�(���#�+^�u/R���W�9�ͮG:F�R��i�r����}���*��Vo��*�N�'�^L`!2{���س�B�غ|x	���m)G�$(!�
��Ł)���/���Eb�1X#y\e^�tc�k��D�.9����(��>��P?n`t0��i�b��|�C�.�,5˵���tl
:{�g&�)�TcI�_�S��.�PƵ�;��'�iI2�:XL"�C��i��9LT;����e��������+X�^ �	�$x��ckd�x��g��}���Os�M�K��Z�4�w4�/Y�9!t$QǠPr��]��C�.�l�2Yj�	Gu�He�rͿ �-?��W�f�u�X���Kg]��?��4����#5��l)z���9'/-ڣy�7����/�D����Y�`I�@�%�4��5��������&=�|	�';.��Oz�w���r5���Ф�o�L8����-�B��Or;0àc����ȍ=�5{������_�V����l7R�G���(�bh�֎��������J���ұ���˹��
od���=Ú���"R"���쀊�������"�||���/����Jg�)q4�g�w��x����<!�����/x���~~���̩u$2h}DK�-.�dx[������`}c�/�d��70�N��y����b��J��J�R���'�w�{���[GC��!�k)'��]n���]�A"sy`k:M����lz������%�uuu%�g�[��Lɔ�Q�=�Cg������Sb����B�Z�^������Ji�j'���^8M)�X���h �Z�!M�O>�^w�j�T��ZW��#{T|�xh�ť^\9����)h���`-d��ȩQ����7i�x��#��Ov xX�W�\���iXN�x{�-�l�n}��E`߬%#0���Y4��I��M��i��)�>�	�)�Z��|�va���#}3�SS����-�N��-��.w���B���Z�!��]��L{�ݹq�5:Ó~��!p��W�h�F·�w�c�q�z��,.�d��L�b鹥[$��!֝s� �J�ly�cβH�(i�F6�1#d�\.��BP?T�ȥ��Aj�|t�,�"S�k�N^��u��&��RV ��=juU!;P�i�`����	�Q���D���˧���W�l��/'���6�;���Z�P�h#�����M�_W?�H/O��x� ���F4F�%��}�\_�V��*5�^�Z�)a��x��-���:v|3��D�����&�(4�a��<c&0��.vYg ����\{��|��u3�R_B�9�Y<}�C����w��z��ގ'�o�-�(����T���o(�5�8T���,����},)�ffԽ�1rd��z{�T{�d�B�״�a��؂�.a�� /�{��#����j;Z�Q�=�j�^බ�9��F�ċC0�8]JVR(8�j�8��d����W�2H��!�+L�o;�5g�V/x�A3��!�D���J+��]���*)�
[�aa��3i��ix�5��
��4���,���e��*�s�0�>���g��Y�cc�u���p�yF��pܹ
�{6Ug$q�N�m��a|F�6l�n��v�|��*4�iO�a\>oCB�r�
�	�����E~�C�DD�f͂s��xV���) �\2���ˈ��x����f�-�^O&�*(,�a1u��"=�AG�&%� �9�9�K:��T��x�f���{Y���LP������:Z|֪"z�&��{�Z�F��T:�����H�o��
p��ƚ�8Ύm�E��bT͓�������]f2�(�L%���a!��-'�;]���6��(���������N�?S��	��������Y(�1�]h��*tW�xs�� �bJ!���Y�Ξ�����J��r�W��q��9${�ȶ$Ӌ�����Fpb�	�p3�!�d3��%ALX�j���p;z���%��*E�)����WgJ�4s_3�Ơ�����ľ�ܐY��� �_�٬��
á�44L|�l��Ĥ;]
v�|m����m,�ޥR�?0n�N�3�W���;���,��E�.�A҆�6�]	�*el��0>���@d�5��u����X&��=���d6�\Z���3�M]SSZHP�i`F�フ�槷9��Z�9^T2�)���P�OC�����-�?�ǘ}�xs���g�C���N�+���-B;C_̑i$;���#9�y��Io���2pM�u/y�Y��ڍr�v��W�-Λ�����,`��s7�>](��.�lw�vE��F���{~���Lj�>�Hb&�L�&&����uqZg�=�����'���>�ֵӑo��eD�O�:{���r�PIs�])�a�!�v���MK�U��ZY��nf��Q��Aec-�S�6�	�/ad+��y�ǣ�����61C����IU�W��u�e�j���hq6@�A�E�6>4�3�E��+�������t�e%�6*��F22�m[*V��o��_�_5Ѽ���DxBU\�/���%-�aY��G%g8_e��������;��ӻ짱.�/���Rs�Z�*�*��֠��.��\���!72����Ð� ���@��@����T"�H.���Z}S��B��m�T�R^�(\C�-( g�Zֶ�T>o�q9|�����}�]-��ΎG�:� � ���P@"�f���$3���̄�꺱o���F��lWU����W�mn��׌?.�3+��8>�{�M�!6�
�V��TCH�y�����q'��۷�O�2#rNy. ��b�IE�mG:Q��F�Y���8�-�&�Ԯ�|�� A�i�X�D�6�J�p�������@u��~�P��o]'BE�>���Ǐ��������A&��;-�N_�X
�O~3)�'֘�觺�ge�_�L��e�ŷ����Eq��:c2��\]�*X򃇅�5/�ȃR"����k���*���� �>���u��_h1�5Bp�d��"��F2�p$�Z�Z�=�N�����ˁ%T�	�L�[��,+ͪ�J]�9��!A��:��+S�O68U����lV9I��'�J����&[���p�Ӯ���t�@��Ј`h,�9�EQ�B��@4���tN�&W���!��I��n͛���rUP�Â��Q�JQj��2i�P���4}��+J�L�.
I�M�j�i��C��*���6�Lq!�l*1����6�3֖5�B*[��"�0>��v����넿����ZL_����_�N�̯��znjG�#��z��>aH�n����������I�WH���U�*$m���װ���Q�=U?픷 ;{ϟ꺺�pS�Od�1�09��X�����Wͳ�9<��E�r�Y�En߀�虰 $5�.I�pE�Q�_�v�G�������冩��ث+P���8��zU�����e���O9�-|�,�d��6{L�(6�4���\�&�Ѧj���]�yz���{��o,UR��r�1�H5���N6�X�8E���X�=�ܬ
�F6OL���{�"R{�¬ҭ�=|����7CUQ���)��"!��B����2g�t��fǢ��Dc�����P���w:v���\X����(u"��h�?��2��'��	�ݡ8�!Hqi�x��V<��/N��B)��wi�����.��u�����uֱ���={ϙ��W�JR���y���$>#�h��n�k�ή���Y^���ɟt�,����k@��.�z����s%h�98L�׊�0�x1nM�ך�����QD,]Ji��N6]�;G�m��
�w5�>њ����if/�͂�p��f��_Y"o����%�C��B<S����YSYx�x�U�2�o���!/܃W�1�W�?D�)�qZ;����YRV���s;*g�=Q��j2c]!ށo�n��e���~ޝ�������݁R5�˘�NuG-y��6W�^[��#��_$�2��J��s�J��^���UD��$��'�[�t�X-G��fa`7����)wU��!�lP��gtX�)� 7�r�?{FԁXY4aS����p�\t��X[,b�@�CA���#�Q�H����.���k�4�w��?p���e^�l�g����(�paC@'�b]����g�?]`��>�˲�.�v�����F����P;'�
����y>��s��[��g=Dhx4�֋�-�>�Ÿ����#s��{L6P�"�@�kxX}[Sht�n�J��{PH=s�O&Ԁo�ݝ��QHf✃5��s[
'S0�=���8F:hwB�a1&"Fa�&hX@dMS+6(�_&���R��Ɏ�"��Rf	����&���bv讶�4��pLK���^\��b@�$������xnh�Z�F��'�&M����GZLDM��L�G&�~Y릍�zz��6�3h��:�_+�[�D����Έ9%���o6=�_k�jU����1_�(N㌵��6C�d����V�@�W��T��)����l�)I�#?%�g���5�ob��I����3~��؋���4�t$��Ee��:���wژ�A��X5��] g��e��^Ξ� oD9���4ữ�>	���gƿ{��M½�N$v�^Mw�QI���w�(�$��8M�_zL�P����J$��v�٤�1uJ�
��,���s��QT3�j���T���;�>�������,�4��~����wԘ�]��]Wk_���9pAk��6��YT=���A���l3���?�Z�)�� 2�kx�D!�}u�������Pj6�Ո���1y��<����4s�VM�;~�z�B�u�{r�8Mk+$�ٸ�ZP̭�6$��vڙ����y�G��]�A�����$$���3�}���XA��Á�FEL�y�A*��_�.���,t�2�v�B����M�Wp�|,�g_����	n�)|�J�Pk*��ct	ǠdA� ��=@�w0��#��g�oOt���l~)ҟ��	����=q[ܺ>~�9��ڄ���P���]%�w��7ћPn5ʾ��!������H�*l[�O�:�3����{_�ѪL�5�P�a���x��v���E��q�֎�EH��G}�N��Ҕ�q' Mň[��S
B��#���S���4)_�H�^{ L�o��䄥r��)���:fK7xHƝ~뼎�6E�}.o�[Ɂ�NU~Tf��uә7+�;p��vA5��i���"��@v��d�3I�i� ��icV�!��X��#Io%���[Xk�HBw�����nBmqL�g|�\��yj%d��wR�=��o_Ҹħ�J�8ˠD���&}Hd �_����ҽϺD�b���v6�Q����ݳ�*�� �<��N�T��W��Y�LQ��S/e�2a	���.��'�����ϣ��
�a"X>�D"�5 �C�kܹ?'cc��m�u
�,���M�̡j�`@��l��3�0eB*�HЃ�y��CЀ����G�J����e�rgH�>u�W[\��8��񍕾>}��Qui�6�x�čF��M��w�g[Ӣg&�`q��t�s7w���K�����Y���>�\�s7�K
���N"�3l;_�|.��KQF�^k{P�L;���Ԕ|:�i�n�1�����J���RGv��i�Ў�R�F{���t�]��M��*���,���{c�!dj^���n5qA�8�|����R_Y+Y��Z'T���Z�H���^'~k.[�vtp��WN�*)����~,WV�cC�~�������
��'��3��
���I�4�ls��\��5�n߿���Ȩ����#3�,s���o�-�H��9�U��DAp��NUFnN蓂A����|R0#��� H�saρ��-z�jY��P��q$𗭭�5!�e�ϟ���44�o���LZ��Z�rGR!�D�	�52**rw��d�`1��ն���*֋I���J[G��6Z�0�n��q5 [$�5��$���C_��V�&i�@����o��m$��&����`f�G�zz�ZnQolzIy�DO�իj�Kx��� F?݅�sI�y�+������A"Qi_�u�P
x����b5r���piT�
66��CR��?�!���<==��E^JkAY*ըC��E�'ǰ�H�Y0�4י��暶 �c䠀�q#jmK6\�q��H�IH:����L���J>$E
�_zP��x���9e�Mh:���v%Da�6 �y92x6�Щ����}UX��.r�a}���x<������32� �d���F��'����k�y�_�`.�{��G��s�|bv�6��N�����B{P������HIyVQK����E�C�G-�i�����]B^�|��Hn���N�$���M؏Ⱥ���J��)/��ۨ�@��;�F�D��}�N@W	z�{��1�n)c]y�V��G�i�à��e-{C��n��[��ig�dĮ#��j�X���ӽ���n�[�@G��-�x�����-���;�Y�-����}H#���� ;y��1���%���X��㏫��f�A�gM$��?���}DSzE���l��vsqV����Z����H��q4]i��h�%۳��Kܹ�!��+�����l5��#w�L�ퟑ�B�j�՘��a���xs�����g,���5܏>�n0p�}����b��ikk�W��$��I��ylR�z����K?��A*E(�2�{�\")���6��L����Y�����܊���;�Ko�*>῱�C~c�CR5�Y|��؍i����t�tdG��X{����8~���M��y]S�B�y�kEz=[�9�ݽ�� 绮�3�5��Ro����e�h���o%��H|�}��U�s�s�n�A�߱,7aR��u+L���wJ{� C�b�z����>�H��w��n�ݯeW��/�rDŘ�[Ź�8�=�\��Be�ȍW?9��R}ji�G{�KM=~6zӂU�K�]�+�61��k9ȸ��[,҅�\ձm�޳eɵ~��5�Q㽘
Nyy���2L&l����Xg&؝�OÇu�:% �`"�К&4؞�v�)4h%���ד�!H���f&[�aV��o(�dUv���Ǻ��Fdy�Z�" �s��5rb9�o4uð���A?���]s�}#�4��j�����{��#�;z��H)+��eۿ�	����?�S��lRx�iCibc�͖�)�3�m���Y�+�q]��7�S����߯t�4���oZ6K�3��I��L�l��=�#&gL�>Z�42������g�9�7��J���sZ$�]�@�9
OE�2^�>d�@8����h����$�~�7~�E��g��Z��yee%��V%?���o;���ֵ��v��y��,����0�1���O�7�XJ���5��4����P��d�#L�[�O��nI�����Hc���%�u~����������H؆M��t*R&;��Ӣ�������COfJ�|��]��!j��Đ%�V}��r� ��<����=��[�U�c�/�۴�8���|S MD������uW�N�X�x*ah�ϙT(��`�Lxv�oZ��Z�:�5B����%|�y�M~&�*��pl��M|��c0�?.=$���Z8�� p㫾��,�Q\��t�ʵy��<$��d���;Q�b�*%[ETꕹ%��+��}�pw爧�I�4�{��e��܇!=�/E8;܏Q�#L7��Q*[�Mc���Q�v�0dt0���3l{Lk�sbš�&���o���g4��0��u�Ry�r��{`�]u��^�rQAI�y�$���õ�*ٌ���O�p��p�w�:�[�DK~�+)�+�f/򾎘�A�T�^F���qQHV_,� &,���#�Q���a�xo�T�Z9$m[�Mz�����?���	�{��R���;�#!�+�C��8�$��ɇ/w��]��e����}�λ�H��Y��k��q�������4NA��V��6/���@�-i_�ƻ3�<P9�b�[M���#&O&��O�ߒ-C���
S�9�����Y�y<9kc����p��6u��9�,�c(hQ b����`��G�8���r:���i�~��.� �i�F�0�>B�QQ�("����o�[���f�#�$rr���SX�vP����)C�-b'%�t]9U�~��'u$�߲t|��0>���+�*��k�����	�|0���̼��Jށ����a4��V
�#�����Q>�)�8�.���R�n"�E�ىڈcs�Ñ�df����l�aJ��?*V����H�_q�d��D�qrrd�izrD�y��S��۲>So�xԈV,����8���>7�NeZb�v���Q�=�EohdDPM�!b �߭�N���$O�ϕf)�䀓���V\eC̍��p����f�* y�V�j�-�p�	�5���G�yS��o�?o6��:-�d��E9L�Ef�Ԭ��p�Td�+4�����+ۂ^��)?�H��ޱE�Ei�ߓ�p�M�`҇������0a7�}�n�)����E����_[� ����߯D�/��ee⫠����^��Q����$�o�2��xR���n:�J��O�G�e�wb���"��R�!���s&'��6"u����F�K���� q���xI�0�P�G���{��m�!?<�׎�\/ 8�e���oOpH�kRDw��#nѥk�Gx�+�C������J/�5�:ͅ�����Np]��=M� S0��DRxיd�2d�lƙ�E�dSi	�A�׻��g����ѥ�r���\��wɿ!bN_����)�pk�47'Ȳy#�����e���X��_r��y�/][�v�֣����᳻���Rx�kG��:���8%'ѓ��P�����Ԙrp`�|6w�4��<��_��n��x�Y�����v&Lil�FN5��u ���L�q����n]DC��et�>{{�h@�4��b�_��;C딞����� %��fg}�ނ$G2��4C�\FC��*@\Z�Fd
b�C	��G~�}�����7�&�-ϖ��[��mq���hI/�Մ6ceo����Zr>3Y7gާzz�(~4FS-�ԥ��u%4Yr0��J�тN�h?���*,�zm�����,��M1�j�-�;�J�7"cl���S��j!c�:!jq�Z9%�Ş%1uA�_׉���TB��8"� f��� JV�#j-@y�>"�z&�}g�o���w*(�(>EwC;�����:T�j[GW�����K�Ϝ���XA�9*�� +�g��գv��(�Em�g.����@FW�CT�����x�h&w�%�YO���Jl�qc��ԭPr����2r���"P�"�eM�P�$�k"vf��!]B��L�����(瓯��h�e�h���.���4*-�u�2�)�4,d�˭p���V��k\d�D�Yx�?���W�^aD0�!�aS�������'`y��2�Xs��u�Z`�q�Uf��~�8}Z��5��(W,G�r���ؘ��<J��4�zV�����z��[�dL����?99=^�o:�c����=�d��!�l4H����F�D<o��.�(>=�7��-܉�u�f/~|�;��7����ەg	UD��a�4ґ׭ �#�� c��2��=�7�>u?v�g����<)�
�GGq�z
�v�$�4���i��,l{��Щ��O�2��Aڗ������K5;;��ם��_۬�%��#A��|�P���]�(�H�~��� �ROȻ�ͽ	��ԯ��V �/���m��fhe ��+\�L�G����{y��[,�$��b'�qm��6
qJo��:��cA|cK�6��d/(�~��+m�L�-�9����l�L��5~O�~wa��2$�.3Yƹt���鍸��M|��.�i{zD{l}N���id��|*���ã
t0�w�mv���=4%��ʉ8�:�j���AV ��/zw�߫�j@%�o��6�<�9K��<��S PaU�QzR3��G���FY���SJ�	"��^e������wƊΉ�O�2�
��CKD��:�Z

�n�9���R�~�0������[��y�L�~ʪ�W˄��Mj[��x�kk.�o�����R�P�����*6G�>�R����Ӆ	�.�c�}I���������2|����X�W�>}�mv2?�/�\oD��Pv�R9_G��/��
i�8��֒�ۜ�=��xVN���Bh��c�_��A�dm1�o��`R\z.�~�D�XH�2�ewݔP��@ã��.�|c``�,�5������mS��ַ���6�����*�A� �Z�⾈bx���)}�J`�؄�T�ơ�m\��ќ`��2���ϋڝ���ȶt�����`�$�����&�{�Y駆 �9��afc���=�`���=���s។&$�|���.y!�N��i���!�DU,��qA��Ч?X��a��}i��,�T?]��>�pG[�B���j���1]����H�M\�˿�Cw��xgˁ�W�<<[#]�8��u� ���绗��o�ㅤ �*hq��oF��-Ǽ�"������#zjv܈6x*]:��|�<�XO6�_
��LK�q��5|l~=���T��s�z�od-�����i�xq�E�i�$�j@��xğ*�%�r���%B��Yj�˸ط"~�$w���mUF��ի�b�",���>�K�o����N�'((�@���T�!�P[���UՌ�-�e����T8�F�U;���r����3˟�Ǽ-�wA*�������.g)3B	�bbbl���|�8)cs1��97pw&/��Q�/4fQ"va�/�w�s">3�ڵX>�C�sy���ߌ�4G�c����{�Mt~ג�Bއ�v��ł��G�B�Csob���kUߝ�2�A6�=vƬ���[�=�2�X!Z�#�0���10}�-�7�W�r���*L�����O2gF��-��1i*�s'h��|<���ZȎ�E9��s?E�����0W��;֢������<JP�0M�v����HJf=���zO�ȭC*I�;!D����|����1�+�d��1�O���/�؂����y��#�t����9N�q�~�!!�wH�5O�>���Y����D�l��O+B>�VF�U�T�{��v~�d}/Խ��f۱h��;j7�ߔ�����ิ�Y���sĆ}���q��,D�����z���x$	]�rö-�04���Ȥ`�.������'G���dgF>1����[�%�Pq3=C$E�y#��nI8f(^p'�W��L%L{�
��&'��o>d�Vp��#opR͂����nÑ�l��k�_�� X�	��;��`�"h`��M�h�S�#<���pV��)��
�Ì��s6FȮ0ʿ�S�JX��~����e��p:�Z��wP��Ҋ
��� 7 ���^�������[R>Yo��ů��!C�cB%k�Uh��̝V�͚�䶀*Kvy��v��������T���:�G��\�O�9;���2�8��`����k} =��e��T3h����r9|���>�(��/=)ÿ�z�Lx��V�j?�������	���uu�PH)��PqA|h���M�&_����G���.����^�koL��{�K�����$�W�"�p�������uur(j���鯛3D~X���{�N�Uo�[���ASY��e�IW�(mz����V�'��9^~˚��GtK|ݓ79r��9n�Ȫ���&_0�/_�0��C}ߩ$��˧Z�;����F���Hf�e=
�}l~�0�N0	ر	X\�۹�9���HϏ��Hz�ݺ��K̃�?5�٦���o�T���e;'{K�}fCƬ�����}�\��ֳ��s,x

F��/�sY��b�zȓ� �;` ���d�M�d�Ļ%V���Oq!<�� 6%��L�{��ګ*֯��#�%Ӵ�qxXcb|Q�W����]Ʉ�cQ�;A���>f���v��Wnl���o/���B�P���q� p᭑�i���H#�
M��^U�Yi�*p����dS	8�^\��T��7�g0	M?��f�R!��M��mٝ�fD^�B��w'(�dd�8��<�����n�����Y�ş �3p�}*�䢪~0S�J�=s��=�/#�Fb8t
��y/I�Q2.ӎ�	��(��>"߻�{��K�_��d�*�C��!?t�7������V[�&�M���8t2�G�8T���on�P�97�-�)���s�L�=�s�������'R�l}0���;1G#�&���H
v�b�P-��,Yi�	������f�P��$R4�}v��XHf�٫N~��Um�g���c���z@�,�÷���	�����/�e �A�=����cҹb����<t �
F�ְ�����NX۷���k>���)����'��&HKdئ��+YE��&�f��('-��(���Y19���M��Ⓑ��z�u/|NK�D�1�+���9Az���t����Q����Uª�k�
�v�-�Bp#jtM��h��r��� �#�>`��қ�mT@T �9��0��b����3�������Z��N9��RJ����F�V�uǄs���9Y/�J���Ct?G��6j�MBL�}c`	`5S�\Rh�W��rNF��?2��uNV�÷���3Q&��z��,O�7�������dz�$��"Y:8p��k{I�VH��iD;��w� ̽�N#�iL]�c� rp�ŗ�SO���0���s�l� ��X��`X�����mb8���ӻ'�s�;�G�#@^��ח�똡��*U�9v(����(y�C#gI�WŃ��т���p���(y��(��Z|����V�
+lv1+�	��ʅۯ��.�e�P�ڑ�K�*�V��>�<��ܩʧP\:�έ�=]U��r��.�cB��uQ~9�"w��p�B^����_T�g����n���6�gӎ��O�����PC'wx���q�v�z&���� ��c�r�qB��#��o�n}w2o4��v�bP��C�e���U�Ce���,@:�2ˏ��C,��՗Dm]
e ˜M^�0�{���r�O���-�녤���7#jg(id��g#��?+��I�Β#������`�i��$��4m"���`�-(�E���4�����~`��l/��b@)mhmD5���� ^8G!<��솷/<��\nƬt�.>G+���%�z*m)����J��h+�7�UVDa��m�Q:�Y,/5��'�_Q��c95E�PS�i������~��Ծ��/���P��@7�KD��+���������J�����­�t=η1��p���<-+��g� �'�댜lT�j鍅|�%wURŝ2���Ha���H2u��H 2d$7� ߊ�.Z��ns'NB�z�IoB��`��k����e���ס������^g"���E�ڃ;���4_THo�����s���g����Nǯ���Twfw�Paf94�ݿ2�_�4D8�&�dz������xw�qF����V�Z*��̼+�$R ?��2Rĝ�����D,��x9Ԋ��Շw"������#_S���a#��QI!������^OI8h ��H�$$͙�r)8xY�P�j3Z�}zާֻ��VG]fo���N�)>����ɩ�������+�(܃S��)]�1_���7�	z&.���hc�����;���ģ��DcMD�U{�|:{��BIމ�^l��-=V�~[Q<5ߗܠ��VDD���r������������F�Ph���fQ�,��ZU�:Yg�]����l��������D���\r�n���I��H�s���ـ,C4�`�x���4x]p�k=�2�91�`���v�,܈/�S��q����(�ңHK.�:��rXDF�&�<z+Vǆ�k��7<߂K����w����W`1x�t��Y�d�R�>S�l/z/m�ѷ�I�ҵ Vh��6���,k����jb._�~ t�Ig�E�~'�3���^���E�:[����f�Jf�e�I��e(��#��ɷ"/L1$?^��SB5,,�$�?F�E��QBwOu�vC�w��@�9�xRҸ)Aȑ�ڷ櫘�o�"l�e�x��"�<�qj�<vL��_Kk�͗��I�;޾�ہ��?{.����W��#�_Z#Š3�uʾ.6����`)�C�����4�{?��mԲ%���Z�D�~�ߐ)?��f��cP�L�S^����3�X�	�.�`U�䃁�4i��u�� ���:�9�'�[����5J��w�������&ߕ����r��~鍧V�S`�]�U��s�I@�l�}�k��"���/d�O��=}�q#¤?a=_�y���.���ʠ�Ps ,S,�������2]P7oj*�5oR�aO ��Q���t�Y�,'��5�"|N�Z�ʂ�����%���B)�����=��O?C�ļ4�ƭԺC���FE�͗U�~($�&u��dy�!��f������*�l(讣h���Y��ˊ�qSmȼ����2c���f�X	��$�9_��ʺ���7���>�w��������h���1���"�&��0�K�U�}>��ҏl�E�Q�C0i䯥�ğ�H�I�Z���.2{Iz��CY2��_��[|���Q���汓�H�\�dM�����&:�~�q�9\j�v��38�@��p�_��v��R�^I���-����2s7���k�m�p��L��C�@����7���4��}�Hݑ��+-a=�2�L�����G-W~��?�s�B�/��g�[�>'γ&������c�z��
t��)��u��{����W����`���OO�Y�i���,���&W����ߪ��b����K���VZ��Y�J�g�0�B�W��c]��k�vA����Ё=K�0�	�z�mZ?���ʘ��c!#�aU٬�1c� �N�c��Zm?��@-��)�̵͌�h9�->�L*��}��ލX3Շ�p���G;%��+M�����L��I��J���2 �W���O���ڵ�������0Sy��^ѽ�;������)u�v�\�3��3���G��P�N'J�Η��N��j�*�եξy���.�X�޳��&��7��{�e;��֛���v���1��ef��v��~FnNL����RZњk=�E��Ed��`�,����G8��`��QE�e������a�jL,�u�m �D��kQ��.�'V�k�E?��bA���>��V����ωY$wJ�3���e1���0���^(D9�ǘ����z���oi�ݝ>�p��g���hZ��zLJ�|���XL#��f�-!S��6��48�����ǟ�U��hJq^`�����:�$Z4
 a=�۱L����i�1l�Hh�+���d�F���R2�ԯ΢�f�][�;Zs�����q�{����kڢ#ɇ���]{�@�=MGA�w�4�0�T��`�B����S����5I!^}_A�+�W|\��2�?JI3��<��İ�c澗F�1OKn{~��wcF�uA8-WK}��/����t�aVo���(����݄31I!����ڲldwo��d��C/ef��ޟ�-��8�����UD���k�/��a`0G�FypK��,sg��bP7X?��9��	�{y��4|R�C����V��	d��(��{\x�H��I���O�|�����оL�+����C�����=���H���G�[�IB"�� ��w�Xt�bu Y�B�=�[fm\�H�>�6��yc���NQC�yQ���`tF�H~�r���q�͇����zz�<���[��qn�1H��P%!Sޱٹ�!d��p%�^��c�y����q.; @k^���%v���e�o������2���ػ�Slv��*���ܥ5.�H�GA��x!T��m��(C\%�\41�6�ͣ�S��A��#��ڵ�F==�N�C�ӟê�[
2����������gR�`�l� p������Ti14(*֜8bP�5��}��`�E��Nh~;J�*y�j5�rcb��%�b�g�Vqo�+�
��K�W���b��hG��U�`h/vA��+��khy[1k^З"U�N"��7����������'�M^��G�m�Ŧ��y��m��"%���<��AOrQث����e_ �4�����9ò��>�P0���Ӄ�=E�#: �;�#�q(�H�z7E��&�7/��I�m:��Fg���\z�tߧ�m�"�O���6��j[�'�F�?z�����}�r�9#�G�'�ؙ�M�;�7577L*��Z�_�<=��`7�k��e�>ˬ���bp�ɚ{�W &��yf4��c�/���|Ku�3�n�⍗v�#��~�|\��:�X��ٴ����\.n�����G��9h��#���6QS�����_�@���d6nF�}ǰ�|�bU�vIj���:~�V|�9;�CK
r�I�x�+g@.�:Z���8�~�2�(��X�M�{���ȹ���k��[(�b<@��6B�:��k�&K����t@Y��P"�E�-���c1�n���z�f�cB(�K;�����Id�5�ώ��MDɲd��p�AݏRR݅���`W��X��a�'���/�տ���~�y�q��w������R�+�6��U/�J,8���r(^��j�9q��
�*Ri����TlCn��._v���{~��z���RV�E:�"�1��]Q����(�a����l;�%�d��ja��A\?t_��F���R�@᎒ƻeLH�#���>2J���ʨ@�6��ˬٷ<E�)����X�[C��;�� �*5m�L��������P9,	��nz!|<��'��m� �d�`ǆ�:	�/ z �Vтt��#:21�6�E	p�l��ig�RUE�Y��6�O��������G���b��@ˀ^����K�����/�p7W�m���c�����v:#���Z��&֗����Q��
�VG�9�c�����M�t���_����@�4|S��Rq��'GaǏ��NwA�?JkD���y�^�c<���GU��p��UI����m�=ɥ�u� !�K�{pv<PX�,����!ϢOmt��'&	4���sC��r��'b��#]�����k�����x�V䡺��b5��]�;�'�T�����y&�ֲu�)榄��7�T�c��Eq@N5 �ʍ������ ݽ��h�L4���FK�����NJ�I�/�e�q�8����ÂҥWd�F� �.b���+t�lW�D׬���a�i�0�d#5��̘\<d~:�G��p��3��}fGP,�ۑh�NS&�9��{@�f�$VLe!���l���;Y[б� %g&`���Է�"�&�z�1�ؗ@g��j6:��7���ҕ�Y��bF�#�H�p��F��h�M���ys�5��Ijg��o�M����17�KEffmI̔t������a�MC��2@S}��p�"������V�����+�MB�;��KAkB�^��Z���EƝ�?�����l�������SL%�5{Ϡ$����$�Q�����W#'H@C��4��_sR��ul�7�N�����B���,:0[Բ�2����u�\�JFX���]9��/�U	�(����/YH_(|���̒� ϗ���.1|��O.�i�_�|�1t����G�_�����~��*�`>� ��d���B8y��I/`� �y�`-O������VZ�4�@�Ҁ�~��s$�Ģe*؉�q�*s�.f�ҡ����bV��E��H;a�%6y��?8x����W�	,4�J(��6�.�6���r{����{5�Y�n�q�u�S��U�J���v���g駏*�W¤�n܃�dg�2^tOu�hP����z����72�z�m�2��J��#�Y��3�}V�} �?r͠��p��7I17����l��:�����*�G$�RM�@i�� $�?b����Eo&�=��w�����o�rT 8��U5s���q?/��M�v!m>;�:��V�CP{h5De�G@H�|v�_�g�N���E-�{h�Uz��ro�ۙY����@;"���R4�_+!����!C>��9��Q����T�N����Z;|��M݋Q�x��Z�T��Ӄ�rd��'+�{ѓ<NV$4�W٢�\�A���LX����)��[��rk�2@.�Ě��&�V_����[���#� /��#�%{�^��|r�ԅ����䴵8��֟���v���}�"C�����0n�� m�� pH���o�(`�i��n�[[��:���aY�I���%;�Y����>,�}���IXh�Va���zq!��t���|!6�����<��7�z�^�OO�X��R�˅��3��|�ܓ�ۯ���������'Cl� $|`�v&]t�L�-]5FBs#���$O�3�-���k��f��@�ze_�24UNtRF��U�xvr�J6�%_����Uv�Z�i ��?Lgw��뭳��)L
.=��N���9�;Ʊ_���� ܠ��*��h�.�4؍��Nk݀�܀]קQ��~{��՟wB�:nі.�YP����Y�����Phe�~q��N������C���Tx��F���O�G�hT����T)H}>�ه����"_*+��a�\��$��aq�m❄Af�V ��z:�uةMľ�'�	�U�Ś�W	B���.�����L�=��2���4;�q`A̼�ۻٲ7����h23l*Z��tl�5�BC)z���J̳{:�xl����B�t�r��8O�e�
N&ы�����?𐽻��4�J�.쵪��^5zR]�EU~{P�}��=��/�*�՟M��#-%
	:3�1�èa,V�݈�'42����u;�tM�HpDƯٙ����Euϻ7X1_'��cP����X�cd���������ݓpBv 8P��}�{N�,/`!�����l���ȌtA(������V|�x��߇�/?0�S*AAq�����6 ��2+��xǾyhj�yd��W�cj?kt$X�l��e���M+S�����i uQ����-;�MY�̛Ih�����K�p��;҅��(�*��K{����9`�y��*�n�a+Oe�5�1�N~|o�H'}Ϸ|�.�ًaek�\&E�����}=��L�BF@V�+گ�
c�a}�]�����V�_��Ƿn!�P|Ұ4��괴1f��\�KŢŭ�V���U���H�!�Zw(|�O��:}:")�)��N� -|��{�n��@���������$�Ϝ�Y kVLbv=j}�����C��y� 8o�z_�+4�;j����7?�����]������
F���PNZ��K��x���^d9u��u#�N��{z ӱ��B$p���M�-�w��2��xMC;��(%�{�o���Z1�EE��������k�@ݛK�D]6R�Œz��	 �pNTfK��z9$�T�g!�ԫ~ؐ�Ʃ�&����SƯ(K+8��Y��Z�'�C����e��fX��J������0��u�����R�v�o?��q귅$�|����c�Ў��w�W5�#~2���[��}�-1��`��Jb���Lk��!�V�"|�,7�k4��9G���W_],�G�l$�ݞ�r��s�������n��޶�����)β��\�5T�,��w���X0� �,�J}�ѕ5�j�m���eB���G�

��9�]��4~�� �Wa���+��>��s��y��sK�`ߕ���ǫ��m�!]`�K섖d��ǟV,���'㖄�io�++�����0��������
M<!a�uX)���/$��䏽]��n8b e����wX�Y1�@-�� �1iLְ�b������*��t�z K�?�R6�����hW9��!������1�>�.z�5Zt�����D�^�h�肨�D5��=�F	�0zo��������߹f�}�Zk��^��u���$�wt�B��Wh�l₣u����� ����T@_t�B��� 7��[cߧ��l���M��y���Y��[4p3
J�w���{D�B����;/����6KI�%h�������Sw9��<]��- ��3�2VC��]C��*���m�F~3v񗅻���3V��o*,�n�'��B1�\�.�o<ݎ�TCY�4��j��4G#Ψ�O>��N3|����U���X6��l��ӣ����	Jc`�.+��P�����T���KX���}�*L�F__$L���ϸ���"
l��v�G���'�����x��1�]6���T	C�O��-�����v�{%���PX�(��_h������7�͏	tX�'S�����8�Y�Gk��a��e4�^q2��Ľț�׀U�^���U�9|,Z���v��&Q��"A��2��t��ҼA��V��r>\p$Cn�e�X��i"eD��㿵�B��h�Y"D�j'�4]�f����*���C�R8�\��%�dp�%��� �ɋp�}����[�I�d��m�ЎE2�$CFJR�*y�֣@c�%s������s8ӓ�^��?JQl&��i�r2��[l�.�燃�D�m�hNt0�1,HNS���5bj���A��xE�);��������/૸/)q7uek�X�8���	U��Wj��`�*�.!� M��� MkTЩ��7p-)��ߪ��c�x����Gv��pj�W*��qհ(��Y�UyɂGK�7���*`;�Lw&M4�.q�S��17�6��r�J14=½�ޝt�* 0��1�3�����H��-�K]��}�A��:���i��`4��d����L��R`�^A�8qs��mn��@& H}�0�vU���zk��aq	$������H�:�
|8Y�]U��rm֥UYE|,u�#{d>�*x"�2Z�㉢��Ș�{hY�������Hy�&�g�o�50�Bk�6_ր��UҖ�$2��H���n�`��6~�)�/N�)W�16�=sQ��B�"N���F�OT$ߥɦ��Bn��s�3�F�r�8C��q�4K��<p6�u������lKIRVf�]���̈��h�\9��?��n�jփO�������i���B�_�=�ʜ���;��a�����t p��У)ʚJ�A�dO��~��R'3u)`�z{��J����U%	��W]Q� m�Ii!KۭG�W)|m�9�Ƞߤ����@�O(�tV��_�I��'�1^H�mWz�H��L�"�h~G"K.O���K۵�)��oO���ކx���T��a�SÌ((��g���!��w}��=�A+���3�����LP.�:u/sIFӂ��*��ᯀ���|�u�
��[��ぜ����${�	�B���Q4	il xd�P24�����M�y�]�<7rO˃�6��
ll�B�}��<��1xn��PCe~�qc������\�M��F(�C�R�x�K��~��P
�J��:]�O��@����?652���D�2���^�Y7lڛ�Q�R?��n�ϗ�a:bN���}=U��|�ܔ�?�9����	��Ei�i�g�#��K���������д�� ��Iv砥�ͽ���D��������������[?w~���ؒ`V�E4��s�|׊k�����8��tѯ_O���R2"�hN�x�?������^��|�c�1�����������3�!�g��%�����������k�"����A�I_�X���������GS�kl��֦Eb���Yj��J�RA$c�K۟5���ϗ��D��[����qk.�cR�������<�}͕%��,԰�$jaJ�6��3�J�Ę���Nx���Ziwb_Z�i�S�C��A��������g�����:��9�({%Q^���Dv�f��=+9@DU"K@�v��GO��_���i����{p��W^:�U���od��d����1�E��k�0	K~x��mإa�)��Z��鍗��
��ӌ��p`"i�"}�U��sS�c<�� K�:���}��ǉ}��M��HCBG��cJ���������d�/����}�7rd@��� �?Ǐ�_��c`���+=�`������� I�dt� ���L�;��C��Ek�,�&9jz�]��$��F���Mj����=�]�AKOG��)���Nl������\��%�����c�V#��oI8�P
�T�[mwV��r�yI�g+]�u��l����\7*q��].E�oV��y�ZQm���XF1'�����V}J�zlW���6J��x��7�φR_��?�D��L��b܋�^��{���k~�d�l��S\�cMS��D�����y���u�Lƍ��>��/q�^tp4NW�1�~Q�h+���D<lT���OH���ʲ�N�W ����?W=�$��[z�����$���q!9-������;5an����O�*�\y���PF#�S�2�f�o))�T���4!��4�BC�n]�R�ab��
�Q�wh�Q�Ju���9S�����/����H����N�t�)�JR�m�Ͼ�C��vs�-"'5/\Y��,�E�B���ҝ	�r£�Yy�ͯ&.?�T3���1���\/�~j�o��
�޲��#mv���.��IDB�tK����'ZW���B!l��4V_S�n4�0h&�&Mr��y��C4
/=�e">�~��͏%��o����	������G+-����އl�~�)�y����2�y��-�fY�E�7��徏�XꂊOg��+�I(�±����l��-�W���I�	��΋��L�Fp��s��#X���G��}�Ji�,U��`����Վ�Po��]���R!�΍� ��+cz,i�X�����@����A6q;�w��hΎ���;Ł�Fݺ_�~��RK(y[��T���O��f�9�w�ŵૄM
G�@���ͳK�Kg6��K��@b�0{
�sy��m�����ɓ��a��g,��d�݅�<K=����3!;�K�Xs��I:�*R�z�zhn�ߣ��%��`9�y�p����|H{�Bh���V��xv��ܘ��:W�f�m�W���s������fh�t�薳���������z��ns�z��F�߁�� �d�=����~������ZE9&짛mS�]�zOZ�B��h3�0V��ѩ�#�{Z�_/֏x8p{~�G��\�aޞ]��`��B0>
��A�Va�t����)p��J`��)�cx�1Y��پ�=���1����9��h _8�y�_ݙv�畴�R�ٌ�CI��G �����^�^0�qBS���٘7�^ؠ��a�kź��#����$��})?I��$L{M��(�޸��ڲ���<NBc�j$:a)�b��p�Dx�ߖ���s.�G��zG#���T!6�%l����(�^��
�"C�1�~�6����y�N ��B;�Hw����_��1�����"��]�[���7���q8PYQe�K�~8�,�j����;�Y@��+��u��Ֆ�7mң�k�d<]����miG��~;i|�r0��5�I<�T�����R�)��Y�t�Jqϫ_��YK)k$��fZ��J>�h�}���9;=��,��a�,#d�`��秽WOy�*����RL�����7��f��xK`*oBӲ\Zoc�`�̂��{Y#�Wʟ>Ț��ԳyU=�ёu�]�P~wN۸}ۥ���F�X��W����>�1�O/$��$��	Y5��o^�����EHx�š��RZ߄�Qꯙ�v���$��r��~vܑr��rM_c���jꦫs\M��/H�`;V�r~�ȋg������Bm�o�I@#�PU����Ro�Հ.�1�/@���)ׂ�S+A�e�����/� �����`eA&�\�4����,�����X��z�o�3������QwZ~MRw�;ٙ� ���%an` �C3x&��5-��ٻ�$N���6i��Ab�C"$F���>꟥h#���(n*�u�Ku�qz.TߴWX>�E��Ϩac�.	{���Uz��=GQX��J���~�|S�a��?�hi` ���y����{���u&o
���ɯ�Ȼt�W^������)4!���H����+�1�g��.��C�f8C��bP:���A�����5J�.���x	Nᝬn�R3���_R% ���%���Y��z
e�0�C�UF���BW�v,!X=�?������r)�o���=�qB�k��#4ip��<ė����>![�Vz h`�*Ձ�s��wZ~�^�Yr@P��g��=�3����)�r�9�~�yO-�q.��t�Dh
��G-����*q}<�E=u3��[���b���<���ԇ�I��m�<��f�]�	��B�P��K!ښ�k�����rwI����l��y�]7yeb���5�4��	�ZTw���������tX#�O�A�����;�=I}��Nenzzd�MkM�R���}�C����qi��I/�C=\��R�/V�����qA�*;<W�Il�s���w�4�x?� }Rڜ�kѤQ�[d�7�3^#�N)4[63U���
�Y#X3�@�\��u���~���vsKv\����z�ҏW�i8�jW�_3�k|��U��{��o�!Axj��b�c��턑�#�������H4�،�vqm�D'��)�I�ˊj?K��p��>7�~�������4�h�r��?��}�'6�ƹ��i����j���c�E��	H����Jln�}yh]�b:��a�]�%�Aa��.���8-!�ϒľ�7=���GS.6(��j����ˑ6�r��?�/��u#���Ө0�@A���6��g�{vh��)O7��w<�e���r���Q�:w�w�T���!K��è�|���\��7o����jtk�������͗�}|��y���~ k$���˖t >���x�0�9{���uM�l��o��̏� �����7��|�Jv�NQsIܒC�s��̬%�W�����!��c����0)�;������e���77l�啨K�����������oi}l3]eC�|s)������������ͱ�w������W���m���OO�����;Ȑ ����m����;���^�����
�PL�Ռ��k@�S*�{Yu��d��v�e��:Ԣ|����[��ML��%���C8�@�󍽁�;s?�*���wY��<�(�\3�i�"D�7�������U��E$����˺��A��I���^�j��p�z8L�]Rh�o��t��� �*֒� ~���} J\���;�^B6'�)��f���u~��&6�j^p.�� H���p�b�zZ�7���0��˄$W���m/�.z�Gh��lvT9�+N�uY?.�f�,ڂ+����OUeIp]�י|�P����y�۶]�[�!���� ���#�y�8v���+��o���:��L���0����~5�Ҍ�.��t$���W�l��`��8�NJ~��3���	�-)��;%E��^$�������Ҥ��gp�Z4-��*U��vݤg��D�T̪����MMH;�r�l������f�r!�Ա��݈P����d�M�`��� ����A¦�?\���aw�[#�b�D>����(��cEMpMm=고}qp�O9���Ĕu��U5�c6�3U	����Y��V޴�� �k�}��%��	Q5r�Gd�N�k�2����L���FW�����N�H�!>���!$#ΐ]g8��/�i��C�Cዬ�����}K��3J�:O} ����NV.�Ïg3}
\�!C�,��L྇���!��#��oA�B��	T%�<#?'>=ȿ�K�L�Z���Oy��EU�����F���˷1"L��$)ҫ�_
(܁��&	��F��r�&��x6�6�OV�OLN� i�������^V��C��>{ �����8w���{A���Y$s55�R)))���PoEM۬�aH�é��J���
At1Ē�Rc��o���0�O|Ϋ�Ǝ6no��x�"���`�
�G*Y�����j֪O6���M,	�c�b5v4��ů�-?I�zK��}����G.r�S���ݴaoA$8yDĥ�ogx���Gz1��ֻ��/f��S���ѩo�LC�[e�/��Rr�"p��o#O�Mܥ�$筽{�kb2�kg7ؐP�"��O������y�������
3�OX�Q��oJ�a���"5mUһx��dҬ��/͕�h����P뺬a�L1D5%0��z�5ϥJ�����˕���=�d�b�vD��!Zݩ��k�pX�I�0r�?�b��� �yG��G�18/U��\1K9�SVW-+��<��B�qt6���SJ�̊f�i����� uOO����M�>�}��+�_�y=U.��zZ�;����/���y/-��H���H��Y)]K�.z�0�j؈��s���5�y�"�Y)4�۹2�=��D"�m��S������~��l�Ε�����Q��G�֨[�0u�қ�Ĳ&H������y�&�]/YS#<0�A��R�D�ի�S�7v6�z_GP	]}Ǜ�sfz�j�:	s�%��u3枫�⿣��=�K9� }!\�I�q0�O,ԛ�w��M$q��r�?#��X�)\V�JA���hQ��e|ʺ�7?��%���+ �P�Е��z�������e���KI�L%͌���g��f�!�V'�̒�iA[u�5y�?D��K����->���0��N��?08�X��:��U�*��K��CM��V���mYn��%�~��c$�z�qKo(�89R��Ų�$�-���L���k�V8A�$V�W�fTq�(�~_���k��H�7���h�}$y�)��?�+��;�GcV�)O�Jް�Av`:l�����C�m��G���Ƕ[и��~`�q�Çy`�C�G�3j��G���E�x͛��دX��Ӽ�	v���23v��ճW�mV��|�*%���/����1��!nvO�1qчDt�i�DB�jL���Ԃ��^cltd�����aG}{u�V�Z���i��*�k65���9�k����\~f��rbbg�O�}��C4E�H�3KԷ��A���rO�a]�}�u�ʏ�Sc�P.��������A�����n�������@A��y���������/S�$;8>�cЄ�V�������G3y�˙L��p�a�@���b�f"��o�����wO�Fp��R�|�����+G��I�g2���9�+ؚq��H�[�ڶ벻�=x�*U��wɢ���Ͽ���̃D�ͭ��?p�40�S�P��G~Q��ɇ��b���899�X�Hu��Ln�X�¬��S�d�{�x�&d��} �A�< ���n����,ԥ��جvqhr%!dA�vXZ��V���n�^���Q��u�M�B���Ю�HW�H�Wu��2K�-LZ���!��ꕝj����9�UL=�N�@��Kիq�F�.\'6���Q�9"���������;Ig�f��SЮ��^�pڭ�׳�!4Ӈ�h�E@���tA?R:0����!�~�ƛ>�``B�����a���Fș�l-��[�C�3i��%�s��u��9����|�L��z�	i�;���yiZN��S���>�-.�1�NmD�˟�>�5-GU�/����UR>����mV��y^�Ƭ%����?���>�2鉕skM�a"�;~c��C_Z*�������k��O\���X�mVJ!����bد�L�~R�����$�R��5'��������W����������!+��#��p����������>��ӝ�0[ҧ+�L�	��ISpɖ3P*x8��J�O�zQK<f�������j��
%o��Ԑ-����d +9a�>p���� ��T-�}q���AP+d�W7I�����&�� 9���hˈx�S'�@��$9�⥢�Շ��>����`��$��%O=�k���o�l�ia�muP���!L�L�;&I�X��c��!&�G
�:���
\��d�wƄ��a���~?��O��1]|]�oN���S���`ZF�m��5f�œ�쀎�6��A�n��dII�}���� F��gL1 _c:7lki�G�J$�FD���C��e�ڈ��1�{��̯p�/(����S��_��$����ɇ�q������_J����:)x����<��w�z�"8b�]����(�g�R�I���x��[Rع��U|t��X��s�F?d�ޥ��X���=u���4e �������	ޣ �?��ò�H�^ؘa��/�S]�,ʅ7�%�Dd����7����t�t,�@�"�$?��E7iM��6V k:�*�N e��.?p�40=���G�!`4�Y��"��Uv_C@xLV{"��������L�縘Q�??Y� ג�Ǹ6~�;k[H	���<D)-�{������;�P��!\*(D]�6"�`s!@#���w,��7���3�%ee��0�����:��l��MF/�u�@^M�UJ�h�|�����=	����\�'y��<R�А�s6Vr�%\:�f��_A�xa���g`�̪�&P.������A���z���ة�kĳbP�w+�����3s]Xa)�����`��&��J58C����1^�X����c�9�s���G�ͥ�AQ@M 1�/��A����=��ILXݯ�v�}�������-^ꆼ5���T;�[�vC`Er�)Q�49t���O��K2t�r������-���>�t��h���K�����W��{��VrR�nD�Q@�?!�����u"�7b�v;���v���"@YF�;#��<�);Ɠ�+o2�c���	�E<\�P�	��(�SϢ��$f'���%��M~�E�L\b�� F�z�"���u�D|�տsW/CR$vݛ�zs�-I�]�2��W�(�fI�G3��X�2�u3�C�<x�xe����Gh)a4��<��d`K��AQ~���雔*3&�zs�����}��f+���?�ZJ��>Ƞ|�йs!�����&'�l'�$������mN��O�Zr���$7�a���r���q[:MIŷ��IO���2Œ�_dBo.���14��0����f/�Oؽ�:��������`����g�2HY~ؾ��R>�:��AN�������Q�p�~�G�_�3��=}&�������@���N�3I��fzY�>h��_��0�_81v�]hJg�����MK�b�����I�R�v5���X��nT�|�-�`م<hnX\�W^Jс���oE�A�'�b_rj��=j�iSqz�*P#��m߆B�C^>��y�L�<�q�����.�׷����z����4,����)��%��q�B�f��I�51m:��jE�W�KM��P	�ca�ߣ-ؿ���L��Y�YH}j(�l�V��xa}�?��|�9��l�����w���|��x�j�7f[ل�r�A@g���Q��#�Q��Qa�H� Mc�?z�L	C-�E�~{|"C �_�Ft��YbkK����_�TdMf���yi�����n��~��B)��:F�8�g�$v�L�p:��
��]�0�9��99H4V���^�����K����A=�Q��O|r��+f9�3�����3H+���8M���~.�
��s���}{�w�3�k��J�s|6��n�{�|�]�ޤ�H�g����A6O���
<�����i�xI�>7����z�c�Sy|$ԮT��)��i'�b�SĆ��aw�t�@f����K��/9�˄-PL.���)ä�<baffF�sJY�'��GwILi�z��sٳ��=��R߾�G� ��L�X����e�'t;������yE��AN�Eֶ���<����1������:�x�g��X��������Jaz�߾%a���խ�m��L�A�$-n�J�M�8�^U��5�3E�3��I}�HP�:�#��<gm�����j���l�ѐf���;�f����?!�Hb�y}8���xе(�V�c�f?|���^<�Ay!�Q��{�����9�F(�G�i�"�n�vy�̌��s�W��W�f?�3=ևG�}�`�!����;�����%ۍQ��7n�I���7n�S4���~����o��O���h�a�����aҡZB�G����l���>�]�a�]��7��|\n������7O��i�j,�[uγ�����:�WU�`3Ke-e.���/�?|2��lAk���H�_?k���6`
�l� �n}�T
v�Z�Į��h�:pX��n��������5?�c�K2��C�en�eS-��*GL\Z>ݞX�}
��5���	4�Ҷhp�_]���� �mxbd�1'�ؾ�xw�x1|�\H/ᅚ(�+��%<TF[�,y�x{�sw�sֻ�p'8")��g�6��j~���=����<��?I�&G��|Va��̋�)2~�oQ|r(���kЉ�>����.������$8cϦ���ƄȜ�(��;$%>4��kf�b�~
X8�!E���Jr��*[�C�D��-<4�;��Z����q_��U��I[k�������j������ m�T���H�����L�=���~�{����s-\�,lSϹv�����d.�d�0s�s���B<�q��AS.��j���|�o}5l8�}��
磨y��?B��^�g�]^l���5�8a6	��P���5W��o�V�r�����[���C��d�~| Tq
�0	�<@0&W\5U$E2�j]�m�
F�xt�0�M__N���^���݇����U⥘S��ѥl�~�m�E�me��TP��V�m���֭o����Ph�
+�[�Y�՞���L�M:��T^�D�ٺ����Cڶ�]�˿7f��hI�ibZI�����˯��,��g��B�ng8���T˞g9oۑD��-��>HRv�����^�Z���f�nw��s�5��LAJ�*
%	����-���"v���e�Jj=P��0��=��e����M�Ne֝�����������.�Su8'��ޚXOe�R���$����a�µݟ��+B�1���m$S���o<c����⯴ő��8`��§�݃��.))�mȞ��1��� �1�+����ؾgOEO��N�~{I��F��^MDGa
Հ��E�\�'��#	���vV��&&�>5���ʓ��'�����>f\/�U�W�N�J�n]g}��Z�s��BM�ͅ�rJX����r��{S������ҟ@�e��K������X6��Kh�
nC�G1:`�~y�<��"�ª��l�'�'s$(�|z���f	�=�4c�<3�����y=q��(�na���Y'U+j�h�^�d�����	�j[D#9�U+'���[��b��˙�ZKd/���'l��x�T/@3���@���f78p�({�G[́حVF��L���t����uǛ�	l��g`7���XfAP(%���L=��m��� � [O�:��h�5����F��	1�s����g(�F3�.2�����g}Š]+\5�r� {E��G]j󖸮��f7�O�P)!�(��8��a@�a�?1n�\�UW��������u�u��궛ٶO������)�B�Օ-��r(yo�Yi�PV3���f�d���VvХ�"����������D�{A+냖'�Z9���^�>9�ؐN#�	�Ǩ!�c��0�q*"[����E�|�$Z�""�>�7,g��=z�/�IrD8��� d2�U�Ɓ�������g��O�4��ߴa7� ����5�7�������#�O���(-�3W��Ky��mm�O��^�{/��<�s˛�@0�$��q�'�R�v�?��+��ρsc����v�p�'~p����?:�˲��p�d���͛>�.�Q�?,>���~��R�.K����f2��}��8��*~r�|2! ����v��P��'Au<Ţj���:M#���?

�LU}�h$�y�ֆ�����fl�_Qc/� #1�-�{,l�����Oe�c;0Y!��/H����d.�e�PB7(��+�N��J%�u��*�7�����®S'��� O�h#v��D>fGq'Qβh��Ch52�x2R�X~��=d���~�M�9P
Z��:Kl�o�gU0-��ٹ�R)�-/Yt�s�xA`�
�!�9��/(��~x�a�D'�˼�>�=�V���m�u�N�6��r�����s�n�6�z���#��C$Jh:�_©�X�m��Q�?�	茗���$*����@�����Q�a�ַ�"�^>�r���P�'�ލ�(�-���컈�1F*W��G'���^bo�ǾW'x�.�/�9�s����bk�q{�����$���BAs�.j�ی�Qzg+o7tC��C��sK��E�?SN���14X�e�1Y�p�J)Ju�$+��p� ��(�+E�UI�-��k|�kw�Qww��N���W����s����Q܄[�Y��Ra)�BY������J�1���sU̍�B���6t7�|�,����|@�>{�=�ep��b� ���W�9w	��4����?��h���z� ��rP�-�z74�Db��m=�#��a|�����̤���!�q��Ӈ��4�*��F%�q�T�c��Փ9����jǞD���Y���ـ҉~y�e�s�n��%�}2���Ϊ"��D�ڮ��s;�EDe�pj���`0�n�5+��0`X���/�i-s�ӒE��d<��3B�%j�ɷ鞳4*���z		�ر5����҉�_��{B��r/A�3f۹���v>�Y��f����@A�` �r�0ђvp�h'-���H�`	W�R�=l�;��۔��=:��[�0OȡԁSށS�$	"̳��r�ԉQЍ�s8��"=� в@jN�a^��V]���\>	B�ba��I�������/�Rů��󙺱���iD�����l��뽴.���;A��i�Q��@�i�k'vE��C�0R9�*+t܁B������a�Lc\�0�N�"�QbiÊ��S���EЮCt�o��A,D;9�\3�xި��t�	�W�L�Q���p� 4"'��*�^�Ռr��a��ɘa�y�����E��\Os�-l�O*��݋><"������6K�7���o.ߨO�e�u/��=ߙ
*�\�v\���U!���N5*����D��&3���Q��v�-v]����*7�G@l�p�����1���t}�*!X��!��`�+#R����wn�W�X�Hf!b|'������z&�@��_Q�ˈ�4��:gw������)�d�ޛmݝ}�+E$Ey�^D�J�y���u���ɤ��LG�����O'�KE�-���#��x@�UT�L��^rs��� �"��Ii�_���1!�4^Ř^7 ���4u�*�5���+p�4��K�g�Y"#r��H�G'�P�hh;1i[M�@9��0�����M���O���|E�ʫ��̈́�{�Ҙ�ϼ!�N0��L'�`@�tQ'�|;J���{�予V���22(l��I�����K��z�ɂ��x�D�waD�H�C�J�<�C5�����𚂼���N���|!	;8��_���t%1~�J�9�|t�x�����vQ	��O$��w��r�ĕz1����ɜkՆ7S�Y1��K?#�p���郈G�>ډ���֌�On�[uI
��w ��o���FI,�EL��0Jj~kT���P1r�p^�Va�W%1����ʒ �-���5ʹ�
����6/	�~�v��%�m�*cy)��^n�S��U ��Tv��ҡ0����Iǋ{���
a9*���S�?��Uql'�\\4һ�)���(�9�(�J��C3���g��?o�W��Z�Ț��0&G�L��� �V(����;m��9�Ġ˙��脣a	�IA��C�}Unse�8Ȣ|p5M��@��\������2��<ݢp�s��H���c�=y *�޾7�3q������u|�8�eR���x��I��?7X�	ߧ�
�C�u�R@�F�����- "��C�Ca߁��.���,@M)؁���ͣ
 ���)�������z��(bՍ�($�[(����A|���u�L����)E�KO���L;gXL���j� �����bHv��xn�^E�|؎I�_�]_gT�#��������=�	�S�CZ����L�!`��K��t�A2Jx��.�Y��>��
����x�#��e�ԯַ>|5�P�x_A�����.��dwE~�� �`3�	G�& `.<�S�E�[]��&�WlA���͞(�B�#��Qy�A��}pa�͆�L�n��=�!/����>T��"s	FuE��?��7v�A
l?��+�#
�3��d˿u���)��@*`�5��Ǟ5�)�����OQ��uv	�xBaoe��?�
*�QG�Mӓ��j�bQ�Z�g�(�w-����9U��}bx����r}KŶ֭���#�~�b	G*e��LC����I���G)+�K�n<Ʉ�ѭе��bU9��4�S؈T�������OF��]4���cDt4�:�\w��Zhx���9�F��wőy񲅕c�{)�a8ߚ�`�^
�LW��<Z e��Y�4�]@4�	�1�#��\Q�YmQu���ŮM ��^*t���WW�!�����8�XLk!]9d���+R��tvR��h��������Mu�Љ���K���}�����a"'q|��g[���#����T@Lsj��pݺ�J�a{%��g���$݁4Y�ڪ��щܽ�UCQ��¼ö��v
/�(�9p��sO�/R�EF�3x��.�
�fF������1B;�]���Q@'H/Lb�d4v�����������tՈ�&M"�Tvc=����ȤZ"6z�[� N R�a9Jg&ټ�a��1�����kd������kTv�ټ���m"�m.QI�V��!��ؽ�=�iQ�N���3��0�f���԰�Ƅ!���\'p�~����b$�r�UY�Dw�~�X�AwmFJɉ�N�osz��̶�����'�+�{�8~�9Y!��:Q+?1!�Y��B-v=�����>�V�f2#�I��.$	&�F�ê��W�:��֍6��K��"gn�w���m��n\�v<x*�:j6-dJt��(KM��=����Y�|�����������c��s�է��bR��@�>b�mi8�;q�,����#���y��#�ce]�yg�a�"a�y�O��T�=ޜ�FYհ�]� xp��g`��]����n��\M���L����i�4��]��$�H�%�)3�/^7֔g%�),��T7K�u���j��p7/�9ͨ�F������&��ч��E�(�cͩ8�Wd7����|�uMp�f�-���?�>R6��Z_�jtDxPWP*����{�sl�Q��}n2կ��5�Np�.waI��`~)s�3��kx)��z�c1q��@�,qV(|�Q�ծ&\�{L��#�f:�GH~8 6���;q�u�,5ScXa㔘	D��%bJe�mL ��T��������G]Xܞ3�X�ǁ;�6,99Uyn�n�$�;kH1�G�%f�x���6B�Y�Y��*8#��h�S{�waCݽM�(��2�9��)����Y���s�nڒ1���Q9qa���g!l%)�΅��{��`H� ��Ivak��W���ǔ�ZI�h�����|�����M��_b]�} ��*��t��9V���*�h=/0w�����Ģ\��u ����(ٶ*-)����N��DD�ms{^=�f�|=�%\DP"s����C(��n��.�zÆ&�}�N�m9�5?�A��$�;P
��A��Ґ�*>r�!e���j#=��Q�:Hp:��8�K={���_]6�`fGj�����!�|�ֽ��a��1'kȷk��s&#0��a����R����:A�q� X��
d���
4oh�������}0W�5����[�����I^1�v����/�2�"܈��X�^�@��&�%�	��_m�=�ݩ�r�x����[	Bx;�z�j��q�'j-qf������X=���0?�W�ͨKe��'�f�/:�1�`'m�L�Y�����G�Kǩ����sc�7��r{>>��ڰ�r,0s��|��(�S�;��Y�$ N��6��>����|��1�*4�3� {��x�枮Ɂ3w"j�N����Q��Tz�gO�0=����>`G���5_�0���"��˙�E�4٢�E���W���3�D���'؅�d����sDֽiOω��d_��\���*�~/L`��c����K�I����Q`�hU|P��2��S�F.�Mը�k��uT���/�#�H����R*%=�t*1t�HI78RRR����H� C��������V����[���Z�5K\��s���گ��}fDE����}��v
T��H��
6����HX����f=�����#[cMx���6.F9a�u�6Y1$�.������J�_���Јx�!9:��D�sb�L�nC�����RO?>%���	�_�XX?g�}�uG�^�P|]+ܺF�C1�h�;��`~�=�l��[�F��	���w<�̚&�KXC�������6�Eɘ�<���p�k���������xg�d��R>qmode��Kʴ $3�۝kYY}B���˿p� imhl�w�ˢ�6Zib�C�qy\�g:���`w&J��BY�ѽa�{;=<f��['$�=�3}�2VD��#�����!��w��%z=[d��%���o�:����RJ�Z��[���0�@m����V�F��'�<W{����C$^'�7�,���t6�I��+B�1Q^�YCyO��[�|o�p�v�Cf����Y{�ъA�>�I�m��7�!\|r��`14������v�:�Ye�X鰰�?��,�:b���:������$�~7�`/-�,/��� ��^_�&M,�$e]�������{�'EF#���7��� ׾�����x��p�
f0��G�
t��� �����?��wQ8	L�>[��^��C����
0�a=����2���F_���ws��f�2��������K��"�����mXa������:n(�9��ǐ�@��R���#��Mx����fbAW�"?P��$����c�h�?Λ0���J\���vnn���,�����N�(ƺ��G
pt�\#�E���p�Fթ��4qc�+��}�ԎZ	��2�Z�7v��h�5�˺(�|z��	�]������$�r&d���	`Ux͏��!�mU��Z�W��4^����I5�������=n|�r�F5����X�W����X��	���������7R�����t�����5Y������6;�����z��K���s_`5w�[����@H�9�i!\#"��vW`0�j���'cnK�%�����*�q��k�P�%��'���τ�_��P�5�+_uo�5M%� K�{�p����0��lq�Xѣwm�k�rOU?�oS�gx�0lf��w�5��`%e�d
��/�F.�eV����S�׶g	�����1��`˺�8eYEE9ϙ�++F���3u:����x^�����kU���Y�D�����չ��c�!�t�wb��T�;�r� @�*��� *ќ	���R�i� ;;H��db;�ˆ����kF�WIy��z�%�{=P��5g��,*�1\�60 {Hǧ��G�@���Z��%
��q{C��LII�{#��q����U���f����h��������Y�{�>���C��3G�i8iv���ƶ�^J:)_�c�,�E�ji�U
(��c6������WR�VY�F
1ʈJC��߯&��2g����$ß��)K�@Ψ[t��B�VRhW�2l�*�g�&/?E���!?	��.!Bw�rH�Ac�����㥟��tS��K��O��ۻ��`�y|쒔��?���/���T����������Ð�L��r��)"��ǲL�Sn(;:,#���h���O���� 2[�i2��zp��\�6���P�/|=�z�"�?�R�&��Y6� �=Q�'p<��Ea�w��-��}9�qs*>��}\�@+K2�\�h4�N�D�B��PVc�w����$ݔ�lj#�w���Fkh`���L��d�i��§��	=!��7)®�i��I���N_?^r;�@+졾o�b�˚W8t'5���Ҷ�5��EOղ� '�f�U�� 1��#�#M&%Ka	tG���n���cd򎨞O�ǫ=̘i�`�j�Z�\��?����-:A��ߩ\����xv.R��8�/ɨ��V4Y�3����zquS�JŶ3JH��]1g� Ȳe臀T�W�4BEvMz�TӅY�"�DX[�ր��o���j�"�_��6�\�����{�8�vT�cYV��.��sS�!crmT/��I�ji)�:<8Z�@��d�Y��4<[/*G#|+�M<�����j�	,nx�v��d8K���R:�UO :��iŵ��@�h���3���T���W結i`h�#[0J
����@��Өl�(�
����%>l:�4V�)D���*�ן���|4�8p�o
U����E�����En����2&().D�Q�ŒeFL�c9G�v3�n���kH�3�5�^f��Ʀ E4�H�l�BI�� (�D��W֑��Kܛ��{��A���Jc,�Tړ���z�9$���y?:��� '�3����@�=@��oI���¬�c��hG��/Ir&��4��;�Z)���m�OZ��
pjiZ��	�'JUbK�_�hz=+����%_�jXk#��,���q�/�����!5��7q����j=uq>��5�����T-�Íٻ�(�.�u�X���x`���o�0p6�C�#���S���_2qߩ��V��bG�e�G���g��-V3�K6$��?H8�I��:%���@7����-���0iVT	��9�����Ѕ5���0����Bܾ��L�T�ّV���4織Z�a�]�_�(�`7���-� �ȍJz��
�D�f�v$G�(Q+�N}�W�́�Y]��bp��@.�s��K�z�^ئ��t�ӑ7��@o���M��b������*ǋ��x/�N�'~4m������[�;m���jLuB��k���/�]�Z{�L�����Ғ%�@AAa��8��������@pvK*`un�קt���q�}qb�	4"��������*�
���t��������hE�����n��%Č�!�ħ=}M�d$Fr�c�lƽ��R��y`I�L\f�uQ����"Q�pV���X�+-�P���Js��K��"�]���"b���A�je~y��8��R�T��D�ᲈ�d^��#f"_}$�7�͓I����)�=Ώ�︵�/ם��:�Q�|��J0���fup��o�r0�!�[�l�Գ SZ�{�}��k�`�>%�^q�x��RG�뢄�<k���+�ɰ'�6��2�,����)�߃�W9o�s8P��`��C�  �BI_�"��C>����5�['�O[3��9��R!��¸�����@!�kX?����-X��h������ކ��g4ΐ: ��\ǩTy/���s�	��+�G��t��ʭ{bdк+7�ސ��޻|��K\@`�~h���aǂ4�q����(�����,�'�lj�p�)*�ʝ�s��g����i����v;�8I[�Ze�� . Zw�?�K�<�Eo����b�(��0�F���&A��&������`��ۖ�|ǭW`��-+=Q5ꈒ>�wm<���i@k�p�R���v�y��	�k�q�;�p⾬�+)�R��;�u�尗{a6f1j~۱���p�h���*�)�n��O����n 䥱�4��tM�zy���(���_�K�cMjjj�K��j��R��yA���<�i���̮W|���9�$��D�
�4� k�%toQ�Gv�-I���s���Z�~�qdד��m|�gl�t�I䇛�!��n�H?1�q: H�\�)[-mP���հ��d|��955����?s���1撞��*�3�P��b�&H���%�#iv�G�_k�W� �e����5e���]�W���%��б�M߲�eY�yZ$�݁N�$B���M)��8�̙ʨ��/���e�80��o!%�ESJK�D�Wn�n�Y��a�b|�����VE�Ju5�t�p���p�������p�C�K�E��m����8�ٕ�7Dw�S% r�A�2���'�G��<Kt[�&��']�u�� v#Z���s�6#�'K�'�тo"��Y��1�ۃ����8���y O@gL/��Vv���~�UtE����;+<�5��k5��x|��0��]꡸��L>,}r�+�G�K ���{�	�"�	�汘�΅������1���7냊����(��I�8�O��|!K�!N�����U��Kf&�4�8J'����$�%'�3��$������_\)-p���%|���h�Y����m�г�Y]���ql	�M��.��Y��y�W�u(,�����\3����n��P����G�0�5�����N[(���7�t��p�of�yw-|��dm�8E�Y��-��s�8@'@l��o8�:
��B����(���g���a�ߴt� }���1����ֽ�KJK�IJ�J�O#h�������h�`kſ@S��?�yt�vN���6w|�B0dt��8rn��`z����Xp9Bȷ��?�w�6�=9)W�#,��n��CR �o�Ž�ɫ���f<d��N317�-	��&dSG����8Rƌ��.u_0g��%�Vo%�����=/��&��	��h�z 3�`��� 0����D_�@��P%8�b"`������w�L�	i�Y�T��x�luŲY��2UhA�^��?��6s��dŀHgb�ڄ�����'8�����I*q'͇2�H��M�ݪF�˩!Afw�@��Bx���/2�����[<I�z��,��wŠguN�ޛ�l��m����Q8v�ި�$�w��P����B����oJ�b/|O��	u�~S Yu3��w�)�Ɩ�E�����u[w���/3�����b�Aܗ:!'�3��ù���+�M��E�!�Ԉ�ȭx2�"�S�bR�Q	��w|,�ڼ��ɐ&qRWE|��"�1=2�[��j&� ����
�RMMd@M�!�j�K&H���)d5���^�$�0f�k�������Ѭb$X��gV)���5r_��] e&�:�릀%�� �Ǟ�F=+{s��_cJ�$~���Y�>}�k(��{
%��12�Xiv��k? ���_�޼�C���z�q�J�D[�z/���Du��(AӀ�>���Z4���;���|lJh;D�$���mwY�NTb��S�,_�t�-��J�"���>��6)+�������>�H�{C��5o�/S�l!�yx4�tёs�>�D.2�#���R���O�vD5��E}��w���e�m��Ϸ��9�۶�Y�$�@}, �'���]Q(qn.P��t\{���'pj��]Q�$҈�ѢU��ia���J�~���;�.ȯ�L;a���4<�����Ġ���b��(�e� z�Q�@��i�<N�x�y���-~K�	�h�n��wJS��/ zK�y~K�g��q�o��1Y�I�b�d}��d�pEŔ��~�[9�gű�|��:4�� ��t������z�C�����<�=��}�:���O���D+�7���m�r?���^9�n:��̋�Պ�ss�ް�s��R�����c]f�m�o��O�' ��8>h���h�M*�����NE������8�&��v�LZ�^鎴mI��I��z�v����7���;*H���et˩O���[���%�z�KA�՜xu�IC6�@����F�l�dUė����v&��C�I:����t>SK��5:A<��#-vy���_�(���%�'h��G�?M.OYD�gSҬ�h�3�s�(�d��Z���̤:�ڬF��y?�|�*a�L�_Srv=e�j�$�z��]�V�e��|Z.�����6�g����tq�4Ҿz#���Uc�M�Ҿ��דUW�'�jַj%p'�W�K�~�O���M�ڛn6gݠj"��_��ޜ?Ou������xp�7���d�+�����zm�1�Iߎ��)�%�l�P)���kw�RXG�+�b�9����zM�����m�/����m�&~Bh9�2e��Ư���;Lm�	�?�x�[-�ǪE���0�R��V��m*�/�+.k�����7c�ڂ��HOB��:��q�S�����,M�B������������(��ο����<�/)�-��UA��
�k��]�[ �����R�q�:���Jx���&�� ��7����%�S�H�q"��/KN��h��޸���Vߜ��໽J��Qpڨ7D���1��6��;h����?v���-jx=��1k�+�f0ͤ-<!�F(�=ާ��C>��b1(���%�����<FN��l/3�[�����iߩ�P}I�3�G/����I�	�3��_�[�Oj_���kiGzA�3���PSN�f�)��G8��w����;���M�u�k0f8V�61��e�5Eى)
�&2��z5�ꜘO�>	��xgtl���L�ޞ�m?���+^rY�3����/=���Q���.;J�M�� KC�^��+�Y���h��0l�hCDvCv�=�Κ�^#ET��5��O4�LQl���҂�N�CE�i9�P��,r�;"�b�, .��BA�[F��Ζ��;�v�H!�Ga7�ƾ�^����O��no�~��)ű�)ֵ����넨�Hi�ѓ�K��T�hL� ν�����s�%��f���b�;2�g�!hh�Gj��4ߌ����|	x�!v�Q���M�@�<ߑ���&�u�oU=���/h=���RUWh�GV���}���HS��d��FD��I�w�Q�7J��� ^l-v�}�)��v������/7'
�mMU;fY>�3ύg��|�7#�'�Ǡ��[0Yw1�i�	A3N�j��_�~�^'�>��'!�Q-1���|ʮ@��Va��^���">�	D���w,o����Dߵ�Ӳ�Rc
�1���H�զc���}Nܵ��R��e�4�S������g`E�UT����}�wņ�w�ˁ��Hq�/�DqT�-'��57�&��-�����x�Kio�n�3�k�#@7TT���>ی��q?����t��D!?5q�M� uAd��r�������Q0xc�xp���у�'�^��b\g�����&"����X?���y�3��mE�,�y�v�ҟ���y��z[Ԙ��s��{ONd���]�/6���<���Z�}�N� E�]�\F�VeL`F�4 ;K�ucrh��(��VF�_��ȫ@�H����;�|��^�#9"�����z��p���63�[O#�G�Qp�����Տr������e�REG�
}�B�TΜ�q�����SV[��̈́�~T�:|Q��X�����6��f�%��ܕ�����iH��]C>0�Ω�C�h=��I恇�(�½��G�b��d{9����o�����:>B�y����,�����4���. yلmm����e�<���{��C�2R#�[6oߪ�����ps��S��MXKR�hה���1���7����n�ɑ,����cZ��Sy��v��z�O�����}���?�>�;j�B�}�h��W*ӊ�O7����<���Ohe�d �& \�?9 �Ÿj�"���V�7�{s�K��gZt^��;{�̆L
��&�*�BX_��$=^/���=��v�����1�L#�^�mBD����f�(�8�ȵpz����N
mJ&MR��d�ClL���<o�i�G�4נ	7�� �v��{/>�~li�e�y��jl7�[1�r����^�ex�O6ypm�D֞�C�m��R���f��-�D0��nVإ��ͺk���Ge�Ƹ��\{G��϶��+�v�nrϽg�Y��"=a��B�Ԛ?^����n��fk �Z�.��X:.��f>�X�	�i�[%h1��[g�#7�h�kפ�6�a0]a,`;sw��������<f��-5��o�:��b/-�p�it�H4��o�쭝��8-��^CQ��RW������ݥT�/��0�깼3�t6�:������6x�ߵ{5(�ɩ��%n���Yĵ�m�'9'~E��}H��:��������ij�6R�nm�=��i)=�#q�'��tT�����������õ�ʘ�UpPɦa�(��:2���`���WI�6/2"�CQ���G��DJ�v���X��*ˏ B-0�{gp轂���[�$uqg]�;�{E�a�$P�9n�IE�"�M����J	wf���ɟi��X"T�nO�S|��率	n �W!]Y�zVET\��ً)s�3�EԖ�[v	b[�F%|M���딀L=K+�N����;|�Y�dǇ� P_Έ�R��U�?wbӦ�=l#Ly����������)�֥|��Q�#�4��K~_SW��:�ӯTR��p�����"34i��Ej�O����BD�z�є���Sj(O@�QȖJ�|��ڡ�X���������CDԡ����W��H����鵗�"����d��m+c�!�2����V�&���p3��B����Ұ��oݸўm�{=ca���4e�Q>O��i�A����cg����F<�ݣ�j�F1�}�J0_��4>�ɔ����~-��b���q�m�����$^��ZN�?�*a�#iEX�3tD�'Jcv����y�s,�	�wu�r!�����7�z��� ��|�u�^�.�ì��q��2��z
t�	I�E�D�sZu�/�����rP���ת3#�}E�MEȄ*�ܐ��w=�A%4w+.��c^�*�9�D�}!̌��v^|�8ɽ��+����#���P�O����?=irQ�#���N<?3Դ�F�ؤ0.��g���O�$Z�ۣYp��s���T7Z�AqU/Ϧ�N&�
�6Go�^#�̷?���v�1Q͕K���J���}$���!������`[C�������7g���]ޝ�Y���o���AR��
5V^4~��((��5��ݲ������$���G��M���Z��r�ǩz./�I�8+o߹����X�A�ˣ"�����
{��&s�����H-�w��*���bгU�2�'TQH�Q*��{��/�j�ݼ��G���ka�����It��睄�blo�"��aJ뚘��i?���_`b��;!d5QqT/���kp�!Q��ke���fp�`A���g�#+�e�Y��7x��y��E���\���Sٴ9�j��+�B]to?����K�dX����vؠ����h�(��KN��ov�P��(��}�f�xQ�DUytu�Ȓ{S:�RD0���[����V����_�ҷ���M9Չ��!`l/�����!
Ul,�nM�)�g�W�y�L?,a���^T3&NpHM��4�V9Ԫ�@�e�lI�(�T��M����y�.�j*F���<oK.fx��R�'�F�d��8i�_:uc֓gM�o���v̴o�*�/,�1�WZ�N���5����$En�d��$�y>íȆ�Ů�R�M&����OA���.�d/e/�F��"E���n�i�gm�N��=����]Ԉ��l�Y�׸��ξ�d��>�!�cmK��D�9r;�n��U�x�Ò"�������U�'S�F�Y3��w._j��Z*�8�p���>�:���}ȼ�����&.h��6�S��	�tN���J��fl�؋,NfyA���F"�	"�W�L�0�6>�����~�)z�4��A��\Y��n#�o�ZϳK����e��=����O9����&w�0h���j	d=��N�`r0߳��*��՟5|\��h�qR�q����~��3��K'H;@�q�73��D23���FE�_p2�I1WK��tw�(��QX����������u��T�YM��^�G/�A����w��i������kZg��4�6s�<[8uҕ*%���F�³���e|�ޛ�"���kSM:Vn�q�Ï�x����V��j/=�셳��ýΊ��50p)c&�ޖz{˷c�Hƣ�la����ZK��mi���'�ģ����W�����<�7D@�'�gU~YV�?0����6�0Z�p\�<6�\�_:�7]��t�<h!�S��X�6�� M�1^NS�R:MpC}�j�j~ܳe7��	�� XO#�s/O�+������@?"v��){Q�?z�B_�빭?��r��(vn��$�6�zybP}��h��j�.����%�*9P�Lr���U݅�ӿ���p�9�J]�jDX�f�7ҥ�[��%���>�OK8�uK+�6��6�^+� �h\#1Qe<��m:�o)�9K�vπoco��X���M�;vH�m�N�a�4�ަ�����NvԱ7y�"�-�lZ�EF]G��>n�j���t?[��,��>EX)��ŷ��	W��B����hUq*^� �|�~���1�qͿ�'l����.�����C#�9m˲/����9�"C&��Q{	��?g�wM���	k�36�f�{��]x�xb@lΩ
�렪��F~f�.��H{�������NQ���箎	24	}���(��z#;�?�v �,*^�Qlն�.��1�o��������t��9�:�4�gU�ݬT[������g?1�[���x�_N��f��8�f��w���1��l�m��x�`��a������Ƹ�@�ˈ"��}P�$����>���{b��;Q ��R�%��
�\�a��AvRS�� �[��
nM�f����5V�"�1!�6|^�}~�:	8������]a 2���~l ;
�!���������覴PP��+Ѵ�[U����7\��?��Wk�r���8���S�_-��#�\ˬ3���Qlm�-)��y�j�U8����k�z&0M^�/�d�R���w�(��V��$v�K���w���8n�C� ɹX�Z����=�N�V���9w��5���v5�G���� �������w�(�!�j�������6��Ewx�^�?��bPK���	��TI��M*!k�!/+�#���n�X��+<�Ԧ{��Fs��&��zD�4$�Ju�r��I~\�1%!�E��)O��n{H����e��RX�K����s�I��5 ��܋�=0л�,N��>���]qg�ҎQ���v�.�ńP��M���A Mk[�W/�m���6`\���Ub�d0\���������c����e�U�틌[���䖰����������s��9did�o.��:u��e������3hN��o�Kq]��*�-2UC�ځ?)��9F��޻�U� _U��òd�j��S�X�J�Yo�g:�Ҧ���)!�	������;����NF�C+`�j��e�k�15��ak��+A�o�g*c���7���Bʈ�&�O=��:}C���9I-��ly��?�.�W�>Z3�B���W
�P���E�^$�FrV��6��)>��)TY��1�4Fi���t�]�N��
s���Sk2s��_�Ao�L�9V���ar�,;�����i>��?����%/�<��e����cN2�o`��|C�Ze����*�c.��
t+^�Q��od�l��0<�l��M,�E��eF.��5|���H�*�m�V�|��<�.�����y����|&)�c�,,���=����Ò����(.a$,�2����[��C�yy&e菓��'cǉڣk��$�vu�����9'R��!�n���(�7�rx�w�Be�a�����K��o�1G�A�ٕD-;��y4h�b����Q�<L�g�L�ɖ:Y�O���X��1���PV$1��
yu{H^[�x�(���z
�3<W�� ��n�<���1�Ī+�1�L�"���;�N�4��q�Q�bz+a����Y�V������ؽQ����<����������(�onR�%5�x'x�dd2���C1���w��&��2����!wg�4�����2>��7k��4��x��yo� ��\��='��:��T�y�4c��1�ĢEm�����O� ~�qp���Țq%o�sm@JEV���� O~�0���`�������SM�q�2����#m� Q��NA��d(���M�a0�D�~��j:ɖ��#�q*���Oq.�b�WL�T�NR��V���@\Xq�Gv�B7�1l�|K8'H<7��ď����xV��-F��`A�Z��2��uS��,1 \کr�������Բ��m�ܩe�鱛���c�Y�*�SO&�����PY����F"y��P��󐺠$ul��+�x����;�W7��9�?�:�r��m=�5 E��4]�o�V��А�1�q3��'9DEbS�ǧ�`ב�*1a���;�\�� s廿}�"3Ð����	=��h9�1Nf��*��D��axH{Y��p0��s���4�p�oծ�h쵛�v8 Z��j��57���p~� ���7���]���j��|ȸe~��i,�W�w�)�Q�]k)����.�����͋��˞�A�/F���Ec��{�mr#�/6��;Ej�Z�į>Ee{E��#��`�_�$��sS�N
��+K���q�K����(C�-�@��%�ځ�s�x	l�wp,{H9R��ŠE��$J?(:�(�6�=��b=���e��H=��d��'�6�a_�/�+ޡ]C�P�Ĝp���i���pif�(��6����$�ec�1�Tu+��}�N����ۜ��=\����b�����=�t�6P"v�e�JqjC�nߜɭ��@1��~	휌o��uG~�b@�LC�YQ�2���T�<�����Y>���}� ���Y-mb\���p��F��B�Oι��6�Oʼ�0��$���5���OX�%���{H�T�'e��l�t�;��T�@��N��V�%�pr�8`cB��nH��W?��kZh�Z�eOd�<g�`м��I���V�UM��ﻙ�Ha����let�I	��w�qu��r��\,R��
�.�k?���y�{%WQ�������ũ�|�s؉u���x�}�5E��'9����T�+�������;�7��q�ܖ��g���mZ:�r������g��?�g|��4�!%6-�����ȧa�$'r�L[1>���@g�h�li�iG�
d��u"p�-���k��b
�7�W)���UL
B;�~�HnҠ/�F,�+<�	~�}���~JQe�7�187�tr�,ZfU�g����#�EW3+L�gl�0$��ur�-�/ik���R�?�p�fT6C�"=c���j���9��~���Sn__���`<+ֺ��\<w�`�aU���r8x[�_�N�Td��0pv��Mt��
��?ؑ9hZ�8l��f9�����&�6=)�gURRRL�~m=6jz:�w`�gh�-''g'�����?��ph��cӱܲ���MM��a���iByߗyA3�~��w��#�9��O���3���x]q������&ݧܶd#
�;�dҸ�C���<a�f�Pysb���[^���N��/���_�I���؋^�?cI]K{���2���GP��a.�\�s�'���0�N�\��a��C��8�(o��D�d/R���|L�jo��?A����X����S��=�����p�i(b�ы�Ix�̙����uݧ8�d�C�I_���݌����"�"�!"��8.�W�q�N��)G�n�����w�&���+W��j��`��e���� -��Fu��Wn%vݘ�e�rծ�.7'�V��b����m�+�:o>�x�~�P���v�c8������L��L%�^�x�8|�0��~K4��EEȕ�-�o����j��%��b��G��挲��bÜ�:�s�1� t�X�I6�l�?�:���X��	�	�L��g��y��Қ��JV7a���/��ݞ��
Y���0�Z�n��n���qu'P��}_x��~>C��Z+K��B�$*b�t�5�	\����F�X?�y2���oo�� 6�Y
�n�O����6�FD�K�Ž�w>���bD��W�U�=��z�N޼��c�:�(0�����/��#-g�ٞ�=�֓��}|%f�o15@��R��E6�0�ے���O2�E9S�P��޷�����v�l=ݴ�E:e�Gy�ٜS�l��.Uf�*��qK�@������"kYJ���OС�	!v��x��fo�+�џ+bo=Nt�Q�n��B�@��*����&�9]W8z��������i��ѱ�����<�R�Ef]f�oA�7eH㖗V$�4Yחy���R���ԋ��&�K��JRQ�7�1���?��<&�p���2Th�V%i�q���,m��c�S�l���M����v���	w�2��w�]��l���PA`V��k��R�� ��W]
���Z32�\�ɺ�M�(�U)#�f�Q�4�2����U���&�*���2�f��>G��}:�yD���[�!������-RQkA{[\d����,��;���t�'%�8�5`z�gqG��B��4&`M�L|\3;%���`�c�m���gn��Ų޿R ��#���SZYxň�* k1lѬ�����D�_�͔9����{�;����૞D�.s��	>^�_���B��5�>ڦ|�!�{U�(�6#�PJ�TM�Ç����ȱ^fi>���[�aghyJ8gtX��vS�%s����?Lo �K���+#��@i"�^���	1����A�	�PÊ2G�Z[���?�_��3$j�����25����*x1L+y���]��31Tv�����%o^f>��元Yʖ�s�N����� D����]K�쿝�w-�_z��}�ё���BP����ϩ��G�ɽD~�9�V[ޗG�}����[g%g!iJ����OGGaLW"�<Afʼ�L���v� �������Kq���ew��-��U���_h��T�U3�2����U���n#4�e�����;��tI):���_CO.ٯ�%�B�a؂�N���j|nm�M�^��>q�/�L��2�4��?�?����.�_i���k�� `��c;ꅲ��P26�:eO��zE��;�|��u��
9��h�� ����K3/0�� >��v �ׁ<
]���̙��K���`��M&��La��������B-����uT`�*LC������R��|��7Ӽ���3z�mƯ7�uG&�.���$C�Tp�K$���R�jb��rc3�������/Q��<�"� sY�
�Mpi_)�b������V�*����1���K���I��>��v��e�T�J�5��>1��NZ�e��Yf03�&�-�/T��X�|[��r�����,�'��lt{G�b\\m�9}Û><Ժ� .���i��!����j��B��I�� �v����ܯz�_��r/�����x���d��a+,���l���}�^�
�����7���7%���鐦�DҠ�īw��W��lt�m�:㣽�P,����'��m����u*twTp2#Γr��{�@o�?ӄ{���@���ީ}y�a3R-�̌�*3+I;���SRlyTK@*�+D���r"���%���f���0����=v;o��m�֟Z���%f9C7}��|1�KYm=-���qF�t��Xr(����^��cn���@�D�T�q�f+ݓRF4BJ� �FHz(�\�1ֿl9�lp��/��S^cD�(�:?������Z)���T��aDw��%S�@�Ұ�1�W�(ũl�7r���L~�ou_
��F@�T'�j�{O�"QK+wv��`RD���LP%VL������~��������oQF�I�/+��K��]�{�:�,������5$6�0#�\Rߋ���e� �c��}�[��U��oe�`��e�%Ɀ�%���ɊYä��K?�Ju�-��xU�i���g�z�S��'�`��s������ �� T:/���y���6���᠂Xٸ�� 5^��`f�1"JzJ��3�XR�kw[ek0?x{���òH`����7�1�D`)OB2ف��R�Av�Fρt�
x-N�:���s�&��5�D�r��I}�}�7L��v��{��RR?�5�X1�t|O��{�1�2���:dp+��X6��8ݔ�U�Q$�y_��,���VV�3��T/������D����������	?:��p��O�]��r�j\M,z�ZX��CF�:O��3Y}V��S�����W���P--�� ,�Um1ߪ'PZo�h�/��v�EcEUR�������7e4�^��p��d��3�q�+#��m�s����>ȳBT�v�b�e�mɌ* `��_�R����gB��Gm�ϐp�%�^�N.�D���g<>r�5��^�B/W61�A�rZ��!�RER�/�L%��y�Z=�s�>u`s^L��	,�RI��L�dM_���AX���PX��9 �U5i�E�D݉���c�X�ئ�f��5O���߮�����C2ր�d/��dF��4�%p��Ap��/pF�~�=��f��H�=���\4&��Y�2�K.�>� ��C��*�������S{��Ӟk�b��@,���-��//��<P�y@ �/HW��y�<l.��(!7�L"l�#~�k��&���JF$0F��
l�MNUjZ���rh���:��ыU 6�w+i��q���窺��-����X�ł��?��{�-vF�hŝd��qA����Z.����VAyZNf�ch�5ZVn��.` �`ND����}��Ӊڂ'(tz5s�o0?�2❻k��6�w"�5K#�+fqV*Y�R���,Aȋ)���0�5��Z�[�@�N�eQ�����N��'���k�SG�hmm�ЛĻ��s��<�����XZ!]�?Y����Ѿ7�{%M"4Uhf���n�m$6�A��D�@ma����	j+HG��Th�^~AE6Ѳ�1 ��qĵr��fc�G���^7�؊�N�s�>��Sj��;���jL
 {0����8��%��5"�B�"k���L��/�SX%MTk՘�'m!2�Q�Vs��MVǂ�%�fɾ�W�� �l�ɡ#��¤�Hu�͒�b�X'k�,=�z�������)�����=T�x22C.<��,�F1�C89���;��!h!>2 �P��y�g"j)/@v��H� a+��v[�m��el\���ꭣ����a�����PJ�c��Qrh�n�A�e��Q�.������������^�5����{_׵������Hxm��5S,���� k���}� ��4��>{]�3�Pqa<lN�;2D >�ᴉ��!9���k���0��e>j>݀�5���$�wU+`*\��t���{�>�vUƣ�2�9<��@M���U�;�"��&�GT}��xh�T���=88����{�nHϙ|#ϝB�!O��C2�"�U���H����O�]�ҧ�g��.!�H2---�G=Bw�Ƙ"s��g�ـi�ve
���1�(�^���%��9Q���.r2=vh5�Q|��Xa흨��a�ǿK�s�J�ߔ��������[�y�|c4���9�/���H% �χ2���խ[������x���#݁0�mw�z:�B�r���94�bIM�Pr��_�)�����yϙ��,��8M�X��.���Q��R�9�U���D��KF`�+�_�

c���	Թ�jKsLj8���O�g��C��[ڠ��KN˾�5z��B�R0���I��P��r);!8��^dүG�������[䜍�D`Azv������8�#Е�s��OE��1��F�5���jD&�.,���}os��w����8.Z/�oRRż�o��f������ �HZ�gG6Wr%�� @7���"�,�L#Tr�Ls6�FԈ-7��r�qs�7���YHz�VL0GV§	�I ��$��!�M����q��I�h*eQ0"���������#j��h���L�*S�#�'*^$��Y�J�l�fc�A;��U�'�*����!/��mi�J$Y�AX�J�&�\
��Q�vs=�e{Z��Ή��^����H�ԥ��b�%d+Jg��m����ۻ�R�0�jvE�ؙ����'{�x��?7`��p�suGXX�mg����X�'[y���
T8\�E������JQ�1�](Wk_�:�b?}�>J�PA
� h*Ϭ�c�2�g�WT@��Ȍ=��_J[�9Z��Չ�/Ap%�Ӂ�K��·�l����Ǽ���n���\�e�=�L�7�(V��4a�OE�>]	F������,^�o�����4����
+�4�!>�F&�'B�j��C?�!),-���2:rbp��-�Y�4�x{	i��E_�5�A��ն�0:�k��w�_7�7?�e���O��L6lr�������c�{<*fz���Z�����Kz��Z����	���� �5!E�,:5N�&L��ݩY��m�2��˂� ���<������.i�M�(�D��7{��w�i��F/�7ܺ��~z�Y{��U����o�Ԁ�R}C�珯'㙁tt���?�P"��g�i��N�����[O���+�[ч�6�8�~���^������5�5�`�5��� ?Ta�(�<T7�����y�Z^[3bi���-0�-z�F�
���TYӾ0Yy���d�r���kZ�}\��;����o�E��un���$�h���=�t���V�wn �����+t�j%M&MF���t�B���a�_����c��n���@��������"�򈋌���R��%byfh�u� �.zd��T�0����<cK�8�wH��+Δ��k��Z�h�����6�ͷ��\�2��{[<�Q�v��>���Q���5�>kaC�G�$�u���S�\gst?5��$��{�s���*�z+2�d1.O~��%�H��&���/��3~�%Q�׆�7.���������� �ݝ�$7��k�!eI]Pj�MQn��q�f��8VD���1�����*IK
�R��U4*g��8bi/�ΗV9Ј�W@���9ڮ'����t}J2U~I����ܘyn�o~a�I�@j�d�d�LlT��/��*o��,�w|�Z��9�8^��e��B�KyK�9)�l�t���]����϶U;X=��4�g}[���t�Hfr��u�4�1�c�Ѩ��2�((h�$t�9a����]VI�\�o̭ ����k�k�ǧ�������[L�2��-S|�R���WZ�H?m�������y��=�>l7�}9�TuU�k���6�n��	繣x���^�GT$�#vQ~h��>>Ьn�ԎgM�@�*f}��7�]&"������)��3���m��S>�����E��P����z�34�:��仆��EWjF`͛\�o��bb��-!���t7�a���_C����"�g�ZU�ΈV�Ԋ�.�H�u��=�l��!��%FŊ/&�,<�T�:Ey����aUI&8K�l�J�x���jv���`4$cim3���5Z�t������3�Q�k�����qA��;��c�;ۚ{�����a�	_M�_�3uLlQH��IO&\Y�?��&3���x�%� �7[n�d� �H��}gj��ǰSkݢg1���̐�|����G1��弦<��CW��j�������n֠Mf����%qA��s�&����#��OB	F���qx�����:y�d�_�<�.H|&?}KC��J�
�����]�P�	%���LH0�����nB�D_Q�Z���8�urz���9��4[���D�:�B!l"n�����vu����)c�����u7��?m�n�@0��;�ce�1sB�IJ�6���.���f=wK�(��F<����Y�/�s|T���@&y=.���⸙�N�o�~~ߒ�R�0�=Қ�J�*��������ST��w_i�!���Ӌ���s!ډFQ�;�����2�t=���nj�������I�����3�V=F|2�����q~��G�d���ܟ��,]�	w.�YDD����\�%d��TAs�h�ơ��?�o��H���u3�QJ�����rГQ*�)����۞k�~�=�~p���h��ԋ� |O�Kd�a�\@)�;��c,��]�8�%S�� $$�`������՗�.�����E��Ii�MY�\�E���li����{mjsN-�c9�GQHt:��M�ip\�Z|8Şf~�hcn���j�QIK	Hׇ7&u�/� ����74��y�*����7C�Z��=Ƨ,J����F�޸�B�Q���W!��&����9g}3	��V�R�Ò���aK	Oo�)Aaǰ�t�0�!`~���Y�x��ߋ=��_����gznG8^�3���+s��3%$�s�_8�ݐ0~N#��v��k��ʴ7�>�t2��t�~�7�&��A��3�a��z���b)v��m3K��������G�Ppf)��k-p	�FagJfJ��>����9�~`3=z<�3?�	�i-����R=�+a~?��������|��_ `)���eR���h��9&*_���d��o\��U�����CR�1H��@ًُMsh��J-կs����X<N��:�{�Y�i���+~�-�?�0Ȯ��2H<+(�J��qV3]����C1��N�K�:�{���o����v����"*�Wu#_׿�����ڝo#�}�VSm(�Ԃ��lٮ��)@���xׇ���v^���|.��	�?_Mp�>}��y��v�Y�)	�.��x� q����^��˸���"���b�@�@�����F?�e* i3�5"��0���;�b=�Kl/�n5���2�j�c�`i��f��$!�����	 �Z��d^.G%��}�ȉ��v<�b�N�1VQ0�?���{\���UR_xUa��R�e!���v��<�8�8G��ι��������umb�}���������f��L�U���C�5o3JBkê���x�M��B\ƈ���������z����(�����h��a^l�O1Ev����~�N���2⑯nRk�U/�e֍�� �gi�,n2�\�" vQ4[]GD̢��1�Ҳ2��E�.28�.��R��S��'V'����Gq�I�Nsi�F|ϫ��c��~��J�D���*SO=�:�~�nZ��R)ʅ��)������|�7��ld���p�!UE/AQ�%p6d�4	W�Q��yF-Q'�)h�U�$��HR"X��+�U�EM'��Os��
Y'Y=�W>�5[}|�������sS��S�fԺ;ت�F����� ]EG����-�����kﲮ�ާ4�eF-�		:@������T������
�D::N�=��{����7*֫��<3��kHo�HVG�{�)t�M5Zf#z��V����W!k�7�E1/���,����u���I�"짟��°Ż;J���+Tr�c��� m5��!�i�q0v��!�IЪ���Y�f'������A?~��8�G�ðq�kF�Sv���^�֖U
�p4�|�6ZƗ�Zg���j�}u�jѦ�P��/_�4K�k�c�?�H]���/(�B1mΒ���[�̓��9W�D�.6�*����d��*E�Ӵ֍��߽}(����R(�x���,�e���x�׎�����O@a�N�������cw�Z>�e'e@�y_�����<��_<���ܣǏ�0?�%��]�=���iG0��L$�6����/�A�QS1�0�?�$�2�QF��^�u�
Yq�v|y:�]W#���ެ�a���#�)�_0i��Z���/�N\'$$psU����:/I�z��h;]�䃥�H��⯴�Iu���h�}������W��WI�#�� z���G�y��^{8�C����-�xĀM\"��J�&��/��>�w>s���d$Y�r�~�����؁��=\�Z�����}r�L����p�i㸙��{|�tp�����r�y�Wܫ�c�v���� �(5�廝�J����1w��=z|�0�Cj�b#�#���q��f�%��;C��
��E%o��b$��oSG��ď�Ձc{M5����+y*��ƴ�C��hяB��	>%����ooƵg�icI��ifFFV��xmjqd�%7��o�HTG��p-f��y�+.�b5�Q���HQp�UZ�{S� 
w^Y����,E`�n�@�����H��C�P� } C�S��^ü���+���}��Ol��K\��|��}�#?���kM�l�[^b�;�Nn���4��S��Au��.��l�:���Ɣ/�^��:xW6��X�FY2��D�ȼ��@�K��rf�r)^<}��,����H�m���7F;�"��S'�B�o�*�u��k��8�]�uG�c��_r#��a�Fnb�Vv��%D�	xI�)
�ku��Q�ZyA�������Ź��R�LȆj];��#N�4U��#!rL
���e5k���%��E��y���Ġ0�&�J�g戶C�<���+����M\j����_�m�]�<�tM^n-�\#"'�ȏ�D>LS�=�	�4��}�%8��%ƫ�U{��lȕ_�+A�*���z�&)�X��2Tt�Ck�?�X�n�KV�������ɝW&��p��z�S�ǳ\������[���"�]��&��
����Ɨa��
��t&[�j˽��96�he�VjI#��m�U��:��	\ht��M��n��4l�&���M�tU#Sk0(k���{�v{�%�wi��%�����6S�^��3�U���[�3+�9Q}I��=1/8�P��\�<��ˤ��C:�2
�{W\�b,�W��Y@w_�B�g��@^%��Ó�^�7��<����/�����J���yO!;�G���P#�:�
ohm�]�|��c�Ԡ*qwJ���Ȑ��,�T�o�u� �6��f���[����{�"��]A�2%d�>��2�		K�Þ��^���g���E�~�/~�]V*V�iڹ�QC�0fev9�5p]#kj��vxM2ߐD�����}Y%S�&�v_������L_����Ս��H��G��0��g��s<��Ɋ��q߀XS���g��T�~��ݵPR�r5�X�ea`�m{�,G2�N>�L|Po0�(/+���d��~����p��{�*�����l���1�{��$�[�$~�'l(��1\��\�#��˦�����5B��f�pk���̦��7e���
�S�(b�<H���M�:S����N��ݠ`o��_谣���l�y��e�d�P<{qf~ZY�
���v�����v֩���n��ד�$��@��V��0�N���G��7Sw�����H��l���|(`��ض�����0Lq!1���c�N^�C���k�tm/)�,L��-�7��9��b ����Ӄ�ܥB�y�����vv�5�Tvd��N�r�9�k�ܡ���Z�U�휳C��#U��b��} ���������fBx�zf����:q%]�@ovܧs�!�j56��Q�_����:b8O�aTxa�`)���� ��r�����:��ֿϴ��Z�k*��"=�")�ǫ���r�������L��!i�$�#E^g�#���	���F��v���~��,s��גA_��`C8���=�e=(��HX����*����
����>�Y�������'՗�fMxn%<Qf�����9=�j���+�,�9닱Rb^��	7�	�|�ȏo9���2��6��� 錂bB�V��L�N��7[�����Ĳ��JA�M&�ۮ�Y��wʷNF$rw��N6~t�N)�0�Ȇ�i�`w_����j���į\2��7�NN�V�fA_D��^��!|�A;`(M�29��0���2��*:>��#�_j�~0�3��^�2�c�f�+�B���Vb���X�#��iI�IO���7J�J#"?�<\�n�<���ؔ�%V`lEZ


xuS����B�ѾC��ɐ�邛_Έ�C$�A��Z�3e��o������������-�V���uxhVOgN�|���;��+��2c�*�)����*�T灺+������\ �u0~� �v���)��=ъ�McTzG��a4}���>*Oe�6vV�2h� �1��+`�<dLfo�����sC=��}�����eZ[W�����t�q��w���y���?�<�s�nQ�)�N^�a��֧���,�S�=hCC-�����R#8�NO��$��n��R2�f�Ah��R�	Nv�&">y����Ѳ����4"`V٥��L�Mb_eٿ�&��p59r! U�lk�.�.L~��=��y���s���<(���̒c�CJ��0���s32��f��"�fK��]?3lv�k�Z׿��9؜*���'f�I� �'��a�YX0��?�_�����)Z�v����¬���9��w�"�݁��s9)u��`���!�_�
����-�i�L1�Tج�O�r����>�r$ח�|j��H2��L���[���U�ſ�dS��T��ByB�LW�E�qt��T�`��_��/3h��$�	������ Ѓ�-���+������ic?�뿝�h�뽠hY��{����(��h�5]���&GÝȿ��I�D�X2�=�^�֯��?����Du=��Vv�/�q��"zrOp���*U�[�8#��j�7��!��~�?���q��"'%�󻫓�`|��Z�Rf������%����0,�l����Ty�>Z����l���`�_����������Ɇ��3���SB�0����#=���MU�No�	A�ϰk��m԰�y�KC���Gf���5�'���D�K텩q[N1�a�XkߛzU!���8�=y�����K�(�P$���� �=�I��Tf���\����˼5򰱴�$�#_w��r��eV�Xه�A�)���+��A�ܨ%g��!jiĨ�w��a{gǭ5c[��׆�1'��EN���#�l��=o��'u��2d �II*o�T��-y_�,��c�Z�?4�[�).��jُ����A/�1����҂�t�7��gJ;5  ��ٙ��{��i-�(�5�p-ջ�EQ��}�?xP���$\h�H����޶�&&���(و�6�w�U#E���o�݊��\Q�#!�Z,��~�R��+����C#x~a-��o����:}}�G�2���df/������|�m^I����.�op�oΘ�2�dO�ٛ�a�g��M=���JZ��l�sBA�������l�'�\��>�a}q̦V_�E�z89�;+��j<-�m��X*�H��ѫEDWK�� ޮ���ԕ�ɋ���,��TɸfrFl[7g�DE=c�^����=��X�W���Ip>*��E�<	K��9;?@�Ŀ��bZ��r �{ X�u�,Zӯװ8nÌ�ˈN�?� ����Lr�������R4u��w>&���UB,�{e���d��W
aF��f�rkK�f�4�m	��E�G��YH�խ8a��JBB�ӡ���(
dޅ�^oǨL}yq�+!�0c(3ŀ��t����D��o.�+�+sۯ}��]��l�#V6�$�`��������1���nr�e[�|�%I Ճة���:����3��x�篤�9>��(>�Cq*��9� �?�����7�F��m�ӭ��@���Of�&�jT}.��Wu��^r٪H4Ȕ���|���L��Q�W���dxI�kM�+������~�Q+6{l�nX?�!�����]61�����&������Y��ŅOx7���a�� 	�W��l��C�	�:�������"4L[��%���ˊ�s��1�I��!"��_�7�ى��}���њ�ۘ�Ik}����Xm�c�+�i)��W���
�8�@P�]Y2�:�,G�k��O
,~6�n��8��NKK��5l�N����~����(^�'^����p�Hr��"�۽����8?�ƺ��?�7�t�a��Ȱ�vnP�e˵�TXE�)9�Z#Lo��x�E���
=
�����?���u�e�յo�z��r��\	21�V�F��üy���%��9��� ց�K�~���j@�w5v4
��V�a�Hj�4���#U�Om`��B�W
ņ��#Ad���:�$R����#�x}ckv�������������ܗv�>?��A��*yA&��p$^3Y�?�(ćۓZO��_� V���9�d�k�E:~������ ^��Y0?tc�R_ q���S�m�?o)w�yg�{?E���m
�|�g���dq
&+��i9��_����!SrLԄ`+��y��qK�?r����6֛d>��o���Յ�Ҍ���X���^ �c^O�$.���e\��GP�tl�Z��È�S<[�ΧjV}�g�U�U+P���㚄����Uny�W��+�n��t��U]Y�a�Bm��"qD�Q"�;^��L�]of���iQr�*+�B4%�s�����J��@�xo>t�O�¾C�_ʔ���eJ/�ϒÞG!�W�SF�Z�b-�<�^��*�@\GjET�M�X`�IN�A �RL�^_�۸x�	c�MD��B'^r�
�(���������O(�Q ��3��-'xj�H�rP`��o��h�7vA]�	C�	Um���N��G~��=�ŧ��Լ�n�q�֯i$�a)�ƈNtܭ����?�*s���Xo~_�fK c�$��*���}Au�L��G�ͧi�z�;ϙ4֥R��,�Y"Rкƶ�T�,��գ������l���F�,���ٛG��y�v-�H��0��XB7��o������j	}0'����e?��O��v��+E�V�
�����@6�ǯ��[��HF����7�.�[<���ƹ�|ߡi�
�arP�y��S$(,��P��[�`J���G�֒��;�����M�G�l\{��Y&p���}���ғe�hɤ�|�㟅R����@���@��`	ʋ�u�<!m���_Ҟ��̓��\n� �����'6�a=���y�m�ð�/��ya�cUjQ[����\}M��a��ɍ3������򬤣1�&==���^,�X@�<Q���K)�e�0��g2��M����"���[�ഴj�w�$h��Uq�f��q}�a�e&�f&�����[Yf�SH�cV�ݚ�rH�eA�9�� $���I��8oS%τ��;�Y!����q�̸Q�fτ��k
I�_�$���"Kѱ�N�7�W'����8Xa��6���#�8D�n��u���
�����-D�gp��;%B��ܛM�9/-��-�-(��lژDUͽ�+����C�E>�
Č՚�$yC�-��V�PW����S�$����{�!h��G�U�K��},��u�4I^�4(!�0� ����,����8!ٺ��8�<2�������G�͑s�T~e�^�� _��cj��(}��ܰx��2uC� x�Tr�șQ2�����?�N���k���&��ϴ�R���W]dY/�u�7J�+@
�I�|�i,��/������*3�Q��:�Wx����9��*|�u
�<ny*�"y�ͧč|h�;R���Y ���o�����b�EaQQ8zzz9���_��Ttx�*����ZTw�Jʈ���Ѿ�5�u��?{M ��^]�����m&=�o�du�m��2����ӹ���а/�j�����՞A�J�2~��0W��4��EMF�zi�p�.�I��vf�|Ba�zĭ��А[z���Kp�9���l����Rt#G��;O�d��T2=�<d���#k��j]6}�Fr���^:���}���#ۨ��҄g�4z)���^}��JJ:%��, V���9J7�~���)����1) 4�>�ۣ�S��X�{/F$�5����E��b(Ag!�
���r���� K#�z�h�,<�4��#k�L�������((���*���(C�ߐ��=A�x$S��Ko(�����K��*��XJ���u7~=S��nCu�#�����Wf�U��~S�&���F����$I�P
"���Ų�^�uM_�:Ӑ^r���2�� �8�D�N�1=��+e�"&�/��^�_9���d&첚��6��Y\,yY��V��gQ#v��(cߦ3��k^9J{,�fHb�〯��6�-"�+�|W�Q�-�\J:�g�[��{��H�5�����z���Jq.0lǅ�� V	�'��%)�������@���2$j�a e*���hVq��������	z��f�ۓ6�qF���3B��j�k��F���MȃW�_r���C]8�����<�=�S R���.��w�=�����/���مNMO����]�SS�?TW�n�2�-��]9�~�YE!ЖR��xu�&:�� �e(��.��������b��b�SJ�K�����f��B5�az��J03|D�Y���H�CI�?@jK�*��$�i�ȟ:�`��WU��r�l���{� ��^e[��E���֫F�J����ðQ�Y=3),8�*+2���Ĵ�Y�� U6�K�Z�>�'[w���,��$������|P������^�#�"��3��x��Rg�{kH0~�z�^Q��D~j�X��
��3���I��9�Y�Y�� �5��~T� �ٯ7M� �x�b+C�ѹ��p�+�����;�t_0T�=�(�����i]OI��%Z�qt�51��@���Nȇ!��1I;=3��q�*ږ��f''���5�h�g���DFV���t�Q��BpLL@+��q˜)39čRɟ�~�b�6��+#N����m�kk��igmz<>H����`��&�} �	�	�7��۲�q��w�$�d�����u�t-8�8�A�W���O�	��z\o�RTF�2
oŸ���3O�����wi��fR�c@c������^������X�����i���w��Y�'.i��b� 2�G��"�:S2[��D�X��lUVI�m��%+>,=�������_�<�09 U�;m�u�d�a�\�ܷ�o��K�O���Д���_����I������Wv>9��k"g��Bk��h9O�3������@����4��B���U�WR�f��J���}ũ��\q
��^w�����ѳ��hG����g���8�	� �JP'�	3�j�+}�4:𵁡E�>��=��4�?���?�K$X�r7d�~�2�l�==�v�IgW��a��y��~K��:��$�[��y1?,jr�x��{�|��%�̨I�r$#7���ϥ��u�I�fb�9+�mh�5��2�j����z��K�)ѕngg7:v�2y����S1��o�2�â��Ga|�)E/�0c@��	5o�(�n-�Ӧ�v�ךĮ7t��D�AŁ��= �β*�B�G��g�X �D�gHp�ך�ԑ�<�d���&u��o�����.4=֞��L�f.�#�����j�!F']gjR�AD�aaEt5h�E!0���7j��d��2�dUt0������{][�j
:#�\J��r��j�|,�[�M"/A�C�4��/�	�������{@�tX�I�%�1L�=�(I�	_ve�FQ�� P蚧p��c"�����.iƍ*u����D���L��Bфh��WF�r�?��Z�'lΐ�Kթ����P����#�gf`���%ۗ�wK�����u�7w7�׻������%d���`l&�e��	�#���B6�k�,7��m�_���|V���T�]lۂK��C��<w�`2S��w��
tj��g6ނ�UU�G�ޝ���-㉭�A�2�?F(Oӂ!�*N��>���ٱ�T��>J�u�!�*V�͙)�)N-�q�|���%��)�V�G�:,A�A�cԹ�'[�H���WB�qxK�\Ѱ�3d�k�'Ԩ5)�����>�t$���,Y�k�_nDr�o��F��+`��|�w�`*�AAK����[cMٺm8)�q�8�Ҷ���c���WЉ����J�%��6�T��a2���T<�{kf@D���P7;��@�i������j��0eĸ����=��Y�9�V� @�5��\6��S")��W�ۂ�t<�rr�R�%T2q�(SVUclÚA>�Fɗ��lCkіog���*���I:����;��֊��o�ڂ�F�PM��B��D�,� |m���3����o}�I��W>0��m8�[jdO��(c�������}%���&S5 ��̓�Yq����Ek;��˼�]�z�<A�G�
���o[�da��!��]�i�������Ul��*]&�عރï�:mҷ+I��g�ZL�ذ�Tr�,X6��w��Bݮ���"��."��?��\ 9�;l� �0r�����-ƞ#_��GD��WW�u��S�ӂ'�l���}�D�|鬤�?c��EЃ�g��O1R����Ux�����k���V7�<���'|�51Q]NM,����I"<3^�?���[st69D��8�U���D�-ի	8|I�(DV�o��%���[���"o-���zR���^ʈ�w��x�S�r��<����F���3Wg��)�#������I,����m��~�h�`@�V���/�iyb�ѯ�Ob��e��{\�
�|p���(�ڑ�/O�A���,��ilLo)V�^<�a8� )}�1�����;[����uQ�d#ꗉ
�q�k<,�5O�p�z��tH@�0�.F���ɜϹ7�/�1L(!cIa��F���^���8�#��<�n�������#�7B�`Ed�^bs=�7n+<|m(�)�������'��o��QU�̥��ʿ)d��WZ�Π7A33��-�ˌYS�+lV�X? FdJ+ѹ,�_77�J����)�O������H��S�I��|6eP��������\{������RL���[ݏ����8�Z�GZ�(�� �dn��	~��T�N�pG��:<���H�K'����q�7>�DȨY��n�S�FB���т�}EkV�����f��^1�Ӹ`kˊ<�����)�c�ƫAu0�x!f��}x{Z������D�B�+HV�:�'���#�V�����Rw��UߌF{���/��\����yD	��������+����S�h�i!M5�������절�
�@�\�B�d�U�΃�Ni^G�Z�`;������6���=J��TNN^G���p-Z�`;M#����)E���Y��4���9�eJ;Q#�.�+��O���L#ą�u�.F��/�����F�`�%��A�t�ۉ�:&K�`�Tun��K�Ss��B����!#D�cR1��&~ ���	���xyX�� �4�!,4ͷL��� V��������lz�p����2ҽ�P�57��3��
Y�;��i��8�"�4�̰U��a)G�_�����:[�x���s���L�gn�?,Ѵ=��K�0�D�5���0� ���*%6��Z�>Sg�Q�s�S�x����%���CG�!/c�jnv�T��ڷX"��C*��R*�F-��z嘖Q��j��\���W�6�z���+r,�c͆t���>Wr��S��b/9������W���e��̷n[�kc�3�ge!�ΉrrrB�E�@�����t�.P�[Ӭjh�g�Ķ��<�[��E;�\�]�3�]$�����mZN�X+ǜZs�a4�JSS�-����o��O��FC�c7ߊ|n/�\�.�nn�I��� 윕�j8A��Xqq�}Yīza��XU�A��*��E���a)�R�3�#�eE5�����%��%1���5�ѕcQ�;zD�N�H���~u��y�}�j���ƀ�m��	�c3�.2���buJ�m0ȩ�M��DB��pX�E
�t�vF:4�o6]��)Z��r�nw�J�RC�^�QT,{¥�g�#�ּ�;`M�ﯩm�����d05`oR9ZS_G磀��8?��4w8vwX��O�1C>����_�s�{��$1Tڢ��W'��#a<����Ү�kʧ=�6+3�q��"��K��X�W���IE��&5&��<?8R���Ob'Whdp�a�|��gpL_�^�iѽ�qw�f�/���e���k�_�c:��mF�#(e�Oj�HC}G���D�i.��_�a<�#VN������D�$��nEx�Nڼ�k�j��|2�g|i�Q������ja�Yٚcq'�خ=5��hG��~`���᜝;겍�KA(� ��o�����U�E��a�Ȥ�;b>��?/��t�Zpۮ���}pL�rY��[A��mИ������������s�Z���w�d���ي����!&�!!!���m��'=5�
�ԥ9hP�l�^a�`����ѱ1t�����V���=A@g������a��wٻH(Y)q������]�L#i,oi[��.��o����'����c���Vݟ��p���s��G�*�6�U��-��%|�a٦��1����Ԋ[��
�ҝM;�O?�P��Q�\*�-��`,����)��y��4$��3@ʍW�1)��J��a*�;�,v�z��7 �Z�Z�,�L:���j:�a�/�;���L�.���eu����Ȱ�����2��&ʕ8�\�� )������q�U�)	o��.�Å�)�5G���A.]���8��l�v�]6�Y�qZlAC�Ut��
#�C�^0�-:����<F=6��We���Y@eԶ�G�^�kO�Y}�d�?Ql��V؝3�C�Y��	�k^��HN��
2UH����ڮ�I%�(��A�}�b9a#q��uH�����*}�L1��q����>����o�`��م�Cm
zQ[y��|/��;R-]�?ow��;��[a>�!?u���</���w�M�g�;�Z���@���0Z'���h�>�\А��3>χ{1�1�eX�'M}]���!���/l�Y���� �E^Iz#�;��/�)����7q�	q�)���u����^���o�����(^s����q��m�{�7-�D�&t{)Ͼ	�i'Y}��&	�xk�nԬ��*T}	.�c�:?��&��y�����״i���M �s���	�q'�p�P'
��p�y�,c�� �)������@䫾Z,�c��ҡ�^���TM:��I��T��Am�88����^��翬�+--��~�X�__�4յ(��o����Ou��9%/�i�7Va���P+�������=��/)�In����;�S�7Sט��c(�lA\���@�f|2�Z��/�zދ�︤p��w�.��R�T����Ë�N5�w��/6V�+����o��ݒ�<��~��Aׁ�wP����rs������IqdNk�n|����"0�پ�+�Kx)C�[�|���^��z<���Z���x���tZM""��NFlm�z�e��q����*�d��t���;N��H�)uEN@���dRO���^�#��L>���9��+��ދ�i��4�����X�20�Yg":iJ2ª�֦E=���������˱�]v?~1�ebV�hZ&K�sۏ|�\�Nd0� �c���>'�([w/��ꞁ�P��,so�㖜�0�>�$�������Z�Z���h�L��aߐ�)Ɲ�9n�2�U�$� �Ҍ�ǁy�`˿N������.[6J�~czf7��Y\C�����VF��S�[]����j�ol�j����.<� ������=[!&�E	
҇;a)L�Z��Š����8�z�(|�7�<����c���X�_`�>_��1��]�W��sQ!�[=��NQw/��qܪo�����?�����{mF���N^$]�.b�B(�|��d	Re�]WY	b-fMz��%���	�E��9��g�x��_����@N�+���&���7���Li��#�Kb#�xe��%/�ϔ�t�p�/��a��G��+k[����/��B������s�8���R<GW�f����c�L���ؖ�#)ɋ�T�X���٩G�e����S�ec�uH��j]SR�$a0�n�AiE����3G�T������3^��S�%ƾ�~&X�46:�n��>bv��0��r��##4<�r���c�-�� k`X�P��W3���A�ZN�B˗NH]������lO+Ÿ$�y���)��c\��-ѻ�E��ܢ��5ga[^f������y�8�5>Y���#^�����L�R��q�"y��I�59&<6ږV�-:8[Z+�Ll~���0���NV�w��m���]/��,Hr�X�_w�&�����n��+I��þUc�~-;"�،*=�^�;(�c;�0X@6�b;�IǄ�'�*�5����=Y�M����'���0�$�F��l]-mT�ˣSR��[�^	��1z4�&��}ё5��	�YV?��~�六�fw��0��IکSΕ��$�����e{�-2\Ӄ��u��b��u��G�����p�u�Yʡ4GЉ5V�N����w�,��q<�]�X��.$����d�~X�؊���B"p�d�+?n����c ,���G��9�����B? i���������s�IBlG���*Mٕo�<t�b�<�OY�?m�N�����~{��jT��?ɉ�D��g�/X��&]��w֥?����4Km+gW,g�r\Ԗ�kt8Z^|�el;zr<��Ц�t�����k}g�y^ɜ�v#��g�~9|-3��H74Zϸ����U�i�zuØ�5I�9,)z���ټ*i�ӷ�z��T��̅H?V��i/����2x�A���N���R#����02�p��'&�uqdt����9�4P������0�>Q{D�����=�𭬇�w�g�KcAK��N�;�w��5=��M܉L�ĝ�� U�������$V������x3&i��ՑW�8���	����u��ڤ�����?_%�,��)�7��i1�h������q��Uw��F�.�Fҗ�i&���p�׏����\YI���H96Z�kEiqi�=��z�2��tXV��ذ��>I۞N?_?ߛ��=Λ�!�d�4j�MVzG�%9A���4��vxfq�lL��X�Ǫ��4[ɫ��ã�<������Ğ������3(5*�CC�?���K�?O6��?�l�4���@_?�l���0�V����6���i�u.�uHe�U!k�3i�nO���ɇС��r���;ꖆ���~
�._���0���+��c ��Hn�EB\��mnlp�H���� sP���������Ǯ�{{p��߰���9�~g9b�79�P ���(���:"���t&�*%0!�WӪW%�_)'^C�d��f<ԷJ���0ϟ�𯁡��C�-��"q�H�j���ʿ�$���El�Ҍ�� ���-;7�Y������s�-b��`3n���K���e`$-��D�ە*43�
��nl��@�[5)�n��$.�mNl��H�0��rd�<G�*��V��X㻲YX�/��b6�q���^ߐ���,c���$ltd�����6ɖ���Qd�G.;� v��*�6��U�`yְ��9~�������;�E~�λI��s��i��F�M�Ύ�J94�aW��Ce�����%ʔ����?JE��Ȗ�<.X؜��mmo;r����;[�L�vvvisc������������@��r\v��(>����VQxlvpȮ
,�I�;2�v�Ľ��:ȍʮ�\�fK行��d�����!:��K�q�������U���"!��_���	�Vfj�4��^��T[E'v��%�������8W�eX��Q�}�l��#�iTy����:W?ךA����|�;��S��j������=I�ʔ�
*��[�Ԁ��GCD�#�	�p)Y�3��֐M��s���]ֹKU^z"�?F\op����_����� *uI4ē]=�XC ���z�#z5?�VW��x�	�����!h֤�ǚ�Wh��1��K�����l�����vk[�蝩��j5�5�7K���MV�^����L�qxxȑ��1�["�`C�4|�*NLp3��V��a�����ck�#yN�9��M�3������A�����6�g*��qC)�2�f�>��r$�<t�&>�zP�c|�&��s�E�&h�d����A�e���]�b����,.r�Xn�-h�;�����D�Y��1{{����[�ؒV,0�+KL�x�/���"�[�L4�$g!�hv��EE�{���^宑M�J�<iѼ�V1�Xh��㏯$�o]�IJ
�Q�[C.�}��c�Hk��!�=��O4�lv|��I�2�f��H�����IԖP���[�+�I�Jss��%��g����4}{�UF���&�'���Y�p%��?�TiM҂����%���~���[��L�A�fAy�@������ 5$��{ppȑ�Ĝ9�E����C��P`d�G�B��@�!������-�j�0#���̉��F�����O������j�">�A{bw9|��UvRՠ���#SE��g��Yce�<b؜���<,p� f9��;�H�uDM�j��������h��������* �0EҺ8kU�RA�9�6/nB�C%�8����Rѡl���	�B�+8-� iU�	ˑ��f�	}9ǋ�[��ЬX�E����[j��)�%�l�Vو�\N50�&��[D�>K�g��"b$�G����#ц�+F\V����oU�.'E_0��y��.��y⎓��9��nin�$���J�r����>H�&h���-�^@x��2������8��m�m�Ͳ�}�T��z�z���=3&c}}�>{�f��,�>�߰��;��,��5�O�"G����,��S����x��4-�zP4ʴC����u�c��.F=�SJ�"��?�����U�Ţ��=�4��h@U�1S����q�֚>SM��Ɂ�?YkZ0�%�p�T��xp~��!F	�W���f�I+xRE�૱LՎ׎;%M=�T��]=S��7J�&��R���y��OU�8ʩ�f���iA���*R���_eh��tl��<����Ț+T ����=l9�
b�@���Ac�����H_[�����R���W�u��Sr�V��I��XǿVs<���b�h;���FWqVW>na>|���[��<؃�h:�LbЄ�I�\s=<��M���hr,dS?���E"�a���;'�X������v�`�ê��"x	�������{�������#�(��^g5{���Q��zT��6oh+�t��g@В�n�.��o��U�V�g��{�Y/���ctY< �\���u�n�z��j�;E��S�2w��9,Zؼ����AՂV���.��� AO�5k��	�v�]�9b��N��;,�ը����y��Y����V��l�s�u�����:�Iw��ݸ�\���
�9D�ё���\�X)�E]m�q�U �C���{�8u��w��tx~�x����է�A�����'^���d���z����w�2��e��.��3�M�0WE,i���CX��A��`rJ؝\�ޅm;;� ��ߍ�V�G���[U�F�U�V�_�-I>�c��P�8�NI�Xt	�2��}�Zn��%Q���]=��;)��.�b@��_763��\Q�2���᯹q>^04�58�Gc�*F	Y7r�V��q(��MBu�n    IEND�B`�PK   ���X�A�>�|  �  /   images/b5136140-2313-458d-a25d-eb2cb312f8ba.pngԼgTSM�/AP@�R�bC*M:����ޥw�^���X�@z�^B' 

H�$�H��f������Yw���~�����̞y�_�y��5Օ�i�ha0����0%;6t�|b���x�y����pzS־�
>�5T�SV慝o��x�Q�W��v���4x\��"x8�<~�Z���������F��$%x���!�����s��g���++�gkO[[7/wok�����G]CoC�G�����6�V����O�Α�/]m�-��]]ܼ����!^C\�::��Yꊡ�&����-��m��W�i���$=m�ĵ(�w:x'u������������ �����111��w�ޅ�#�^nޖ�p7����_�<����t|��������r��r�c����C�����Kn^�]�@��;���w�P�Ч⚎��.F]���ߐ�')�����㙆���=���癆��g�y�zʻ������gf�;�������m$����,M+)��L��5��US~ �럲<ES5˱���}N��e��s�,ݬ�}�����R����O�f�G�7B�����xo����|���"*xQ2�J��)nzA��O+��$;�F|��1��j�OAa��-r���Zkc�[1���n�M��v���3�4n9�h��"�
u?9m-w�k��{�K�X���__NK�u���v2�!�;nSI޿�v(�6��%�|������_Be��H��E�zt�۷'�:y�d��\�P.�i����Y��[țr����=F����1�>>�ɚ�l΅��}���������%�z�J~�z�O7[��/��}�cm�gR�] ,�BՒ���.�<��Y�[�K��<ezx��j%�<��5
Al�����T�!ye���٪�L� m���gjL��=6�o��b�m����j�SO�Я�#o��<=V��a�y��E�+ļ��\W���i��Bf��TC�r�8��CK9������o�AM�N�N��������c�*��Ȁ�c�Rhz��������dfN��
=\��m]��f­�;���O���i�k�������h��p�	�ix��>���S4ߛpA�ݳ��]	���w7��:������6�*
n���U&By�X���E�q��f�F:Ǹ�r��tiGV|Lb���+tqs;��;~���Hk�8'��ԙ\[�K�#o�!V��w̼��GJ�$�n0���А��!H��t�Y�:}?-��	�*��z �	��?B�WG4�y�A����
J��Rļ*H�I�N8L��ޕ�m�.��;�;x��/�w�G8�&\kХf����а�$p��3x�jŁ����ПU,����+�i�Ϣ�!���J���Rqe�_
A�n���*]�x���膕��4Ɉ��bG��L�f�R5Ⱥ����ࢇLl;#�F3v[��Dry�v��x������^S}� ^�|8�m���`Qe�V�J��y�=\�2���R�7VlTy70��Dfڬ�t>�o�f2�w�[t"���mP���36f{�CC_��ܤ�ʴ(�%�ς�gH�*�l��wXϠ.�@��Y����7f3�7t�3��Ӻ�%���+{�]'�E�&�-�e��j�P⾿�Z�G�f�j/�K[4*2�.��7ɔM�!և8=���4�d���R]r�AW\
5Fb��j���Iz}��_���3��O����w�TG�A�y���U��f�;���*�����*q���I��T����U�rwg��,J>�u�j�K������!s�,;�陻h�_l$x4XȌ�����r��x���a<
;�Q/�t�7W�"G�+ڝ,�*1�c*���������~�
=[���RP���<,����Q�%r@�2jm�Ԯ�IsW�x����M��F�lrGɵ�®�!脌3*�e��i"^~���#����Y��:�M��7��.��d�!��~��l��X����ʥs;&�Mq���y�qZJ�qã�ZDQ{�����^s=�g*^t�9B�W��v �̸�$�k�a���xg��ӥ�	?8�[��B�4��뫳G(�6%Z�6��e��M��3(��ѐ����'�^^�2]�fO�0_N�������љm��Jvǈ-�i��|\��������1^�u@�#�ZNY�Kh?��{�;W�(�N���e��$v��u������v�H1)ht�'�2z;�&=�&͞�]?�ݣ���R]�75GK�T�%����A;���������V���4�ѿy�x��C����K����_"�y�2�Y����w ��Cmx��4�C�����/Cm&�&߿k�2>DGR�r̓�[VÑg���Њ��������(|�4a�n��q�gǍt��I�T�e��I�4봠<q��n� -���7��G����e��;u���|_���gqHy! XP���E�MU�Q �:��+l�&]���ʩ��jm+�؄��v_�
�`gf��T�w���(��W�}�G���^L���V�u�J�y�rǺ} ������<ji�Ȟ]ܻ������ww�t�Z�5~z6!��}��#�J�ծP�E\�]�+r %���)3��4{�@�2=�������ǣ��nk�T@m��"�� ��X<�~C�q�����;̡����C�3*�������3
�K�{%K-��8ò���.-�U_��w�`_����Өm3	�Sʷ��*!�	�=�`��ϗ�g-n�zk��X�H�7m�H��cr�F�d��A�`���u�6@誃��1 �������տߔ�>���з��l�P��y���3��J�x��Ą{���h)��z ���Oǿ:6���G�]eU	�R��UL�RLu�wҘu��m5��)����Y��c�)-CJF	5e&������J�m@�ԩ����q�1c����X��Q��Gˈ�CȚ�CdᮄGm=)p�8�;o�@ �O�Q�*\�S�e�Jh��޼�~[8�-�`�\�Γ��J�9~��M44��{����G0��[�]�k�P��t�*�j�����vW\l�W����;*��K�#��Q'8����^��$��=Q����{_�����mT�T;��-ТF��󨷴H����q|�	܄��?y��a��]�z��jv�(��g׷#�T����Ņ:��j�`�i��|�����ݥ�`����Rٻ ����>��L�Rݧl�F������h���а�'��6+~���^��>!wn�d�a9I�t��g���@@�B�ϯ!�c�V��	��J�^z7N*�,�`�	�xˍ��.e� �G�//^Q>��)
Ҹ�l��-O�>d��(�D	قj�y��8'O��*`V/T�<\b"*h�\k�)�F�n��Q�g�¸�H7֥�4�8���_;�Ǚ���S��H�գ�g��kd�w'�Y}D���)�~L(����_
 >��: �0�r�j���a�1�������dag��	6qq��ya�s�ү�9[���E�+m �@p���4��{��Ɏ.2�A�� "��D������.z�Ps:��Q�U�U�WK�ѝ�A������Ԙ�:�׶��	;ٸb��|��6�Vd�����h�������쒋�y����b� 3�i�A��,��}��L˷es;��|��j;;�y�g���N�)����u��xU�Cs�%��}ru��Nr�g7�a;G褥*��ș�i��LIiQQ� <P��XL�Zr|����Q�(Z�lC�?���r�A��T}5��q�W�V1��T���{7�}�
����Z�^�����#rtx-~-1���
�l�G��+G�f~����C����d�02b�cHKi<�A���뗗1.-�ߢG3�OPƊ��Ԏ��N��"��������9��ݎ伭�&9���T���E/����g��:hn�<�i��>||���L'���]��D"�jP���;nڸ�����5lB߷���~r� �A��?q��S��h�����^^��W�ear�%M���d��Y��o2�o��
=�P$�˓	 ��`dH $lLa���7A�B���-+����\����uS���!G�@C�́�]$�5�sq�4�ҩ���*{Z!���Y�7�zR�e���~������ g�K�yR_�j��[y����e�����o�A����-�H<�Gj TO���s��u����:����z����?�[�W��z��!��7M�,�A���Zcl�>U�ֻ��F����`���v�y���RS�	����4�Ӿ��_�9��g>�S��/16zǭV�K��Lf)D���ǃ��N������M��q��-}�R�f�m
����X�� �5�q;(�0�����ּ�C-�Ͼ�>��0�d�*�EH����/2U����S
·�x����ژT�F�b(��䬿E�t� ^w���X� ႃ��`��G��m���:P�[-�ƺ=����A���3R�{��T���.�f��H�<~Qv�!��iࣣ�����t'�w�ýj�� {�X-Y�������~\�D�Wb�$�3T�P��P��)�ۙ�<�i��k!�z��2N��ͯ!� ?�p�����Y�-�c�Fk\�aܴ���-C|4x3/`�u����X���R���҄�	vWtܱ���dt��;_��n@�>���7\�纵8�RiF�h�Ɓ��B��]`X��B4,W�D���[�0+W�|�nw��Mf��՘*�9b|eK#&��Ã��Y7��z����D�n50��M��eC�|�#Kj{�+�AH�yo����:��앴�$���l��* �d��~l��L�e.��jP�S����£�3��l��\�7q�Ab�Jz�F�wG]��}>S1��	�<�o��y;[j�ȁ��U5��q[X�:�h�E� �����/�t+~5��v�B���W�q� �I]�h��r��n�yj�KO��/��Ѳ��^���S�2������Q�$����ao�y2q�x;���4��}$�ٓ\��Da!�锖0�ӌf�A�C�h4Rp�<p��)ֻ_����$��42��7iJM߹g���gd�j��n���|�y��v��}v�$�y������C�²r�A�k8/�����,�VҼz�V����b
\_�<��N������� �j�|'�a��OK�<���IJIR���+C ÚW���A��Ȇ8�1��D�����b���ԔB�Q����� $Xy �p?��XC���J/k�$G5���_��Ȅ�`�^SF�|襠���}9Z�s��$mmo5�DѨj�7v��o�����	lx}oh8%�gǍ��j(`WC܁C)2({��s�=_im��Ƿ��^/�8�����i��v��?�^�K���o
��Sx�@��H�>N[��/5׬׵5�
����\�[p=]��`SZ��7.�wxP��h�� x���~K%5���tf�����j+��+�� 8?��9|{�V_��zH�rd����|�@��&�� �ԎS�����w5m��_�V�`gF�{�L�jm�T�-U�����|e�����4�CtN+�_s�������Tz���v~EL���sk��-�D�$'T�i���~_XD�2��o1�ث����	u����i��O:o�A����9�N��(6	7���7^������]�N���6n��,ρ0��{L�^�%��'?���8�U�۹����Ru؛|x��˅#u��U�4�[�*2�,�wZ������'X�ʅZp`t��-���;������$�b�Y��+��'�e�p���KO�����z���K�q��R+Sƃ~��rQ�'-�7��ӐN��s���'�b��o~������㲣�;�O����q�k6'�����b�Rhǆh�� �6�AD�/���*��o�q)L�;E����=�wq2׬rp�M5��Ǿ%j�~��ar��|��̾q��έ����e!�'! 5}D�;O�zS�`�]���Q���w\��6��$��7��xPMT�W�1�8W%0:�=�Gj���X,�;�#��h�����s��q����t��n`
���+���`��5�����(ҸX =m�"�y���RY��`3FhM�n.������w��7��f>XG����Os}xVE[}\���-ٿ\BZ+��(Hɱ�u0ЌϞ�!�͇��ɠ}BB�V�:{M�#��3�bcX����G<�[��u/��^i�>$7́�J�	0���y����O}�90�鷌��/�{��(�Ny�^�g�mW���ZZ�2�L%m��~��d��
t )ͤڅ��g �D�`i��!�8��/F���f�; �i/	BջYc�2*iX���gG���/�nK'�; �~���n�������e�l��\!��x��!VƝ��Yf��ﴶ�����v�QsX��w�k�L7�� ��A���Aa1��'��̋�z��B֧��PiGH(lQ^�j�8��ϛ��|!+��>�	(xŪ��Ѝ����񓁽���:,6��iR����Nf�	��8� ��N�IK��ϴ�qi.aKA{>��f�٩��4��]I��V���=�ݯ$�� %,ÐIOgRmt6nî����'@�&�<9����$�r�v�Q�s�!UTO"�Ď�j�jO�Rc F��$�o�V�s�z���{�i�"h}.#C�8[�C�����X�n.6͵��ݭcKUKv���ц5���H��a�~��	`N�O2�w׻̒��&�y�n���i���K*���Gϛ.�`�ⴼ���<P�g���}
K�D�+����� ui��W�Zh�U)��Tҿ��z��b�Ow�;����4�%���H1_���%<����5�#����%��5sN�U���s���3�� }�'@�T
��>�ى�0�r�)���: iND�Q���*��ջ$VZH�=�L���z�/�濞=�w�� �6�f�	^s=h��kl�B�߅	>C�t�@�{��!�U+�{�ܢN�l�|B��_���ְxW��o���)�Ĉm��LPb x�ಊ�\ݯxQa�m��Ѓ�i�������v�y�[�!Ի�U���o��~��s����ծ��ް����a�����AD/pbқ�(f/����񮘖�	����][a0Zep����ʢ%$��G�=% tWP�IS�)�>CZn�W}yA�4F<���eq�)�j�����B9���%|]�&�����
-��Ż����~��=�����߻�2%���c)W�T�r��0���bO��P�-B���N8_�I�����2W����D�݅���04��Zي�^يQ�N���W�����m�֠9hk�eb�^�q�ke Q|��N�!��X6�@�"Y1����2 �ӒyF�z�j�:C)p�M6Њ��G��Oχ;WWMov��=}��Q#]z�%O.���F:��Z/�X`D��-A����8��=�&:�>�m��Ԗ.^�)���I��%��N����4E�6���_�|H{�1��X[�1J�k[���'�@�~�7������h��Myv
ɻ܇v6 f,�x�x \+�jT�zėnw��k�
��8���]2ު΋6D�q����ݜ��G~�Iʂ{3���!���B+bF���U��A�$�}���.��|K�O�y�gڈ3@��@���"Vo�v�ܰu�*k>p��F㜰s^�iE�7�g�c�>�`�lwj0'䓝
�Yi,�@S���&�|�����q�}��L�E���-G������C:�;�f��/�ý��B"$q�o�vs�"l�\葹�,k�nBb7f&"��M���y�8� ��6v4��h��i��B�?J�1ͤ�D��2��{�g�P;M���`ZXi �����-�X{�w�$--����PӶ�enT�ۜ� ���L���w)2H���i�`�u:�oȝ��
��ȡ�p��3�LOв��|S�]�{��x�[����x�L#�3�)��9=�\�RG�������z����%`�ЀCXc�6�8�X=O��:N������M��E��*Ĕ�����yiN�����o��؇ׇm� �V#��@m}��M�*�F<jS����H^?�v<�jp5�^kXeyml�[Ay޹���~+˩��|vn}N3=�y,)W-�^.�İ�R�̕/Wd|r'��ݡ %�,F�A[��\�p�������(���o&���{�ڋ��|Y�+:��hP���d����F��b�Y��t�����*?C���h�$׾�7���5\I�t��W�6���Ik�6�ă}��kF/)ޅ��H�V:mRoO������z��G��*")$��R(Onbܳ�?��o:o^V&��dJ�+��D�L��(��;e2}�pq�|�H��_�i��mr�'�7��.� wX�҈��#�0���gA$؉�x/�Q�k~ĲnU��r2���	���F�a-r������@�Z�L�=�j/��۰n�ྈ}ϥm�SJ�Z�A�b/m�=�=dq�8xn���#At������1Q_��>6�U�ͺC%�\�e��87X�4f�Pc�(��\�9=��6�&�a�������%kT�vhʪ�\�mNí���Y�[���ͦ��B�@��$��,���X2 �����p�UQ���|��EN�`g�/���d�L,=�	��ڙ�آx[��;��i�4t�oZjy�[.90W��X4u���:�!?��oC�̻�s��
:��#5d�g[�P�u����wj3�=c�j�n�-V��3}�џ�)2�p��n���K	m&k�sY�<U#���bd<�Y�MTKq�f�"�����ą��σ�t�������2藜AcM��i�����yr{b$V��|T�j��q��I�� �E24��@�*�k��ݯ`�h�O��-/ln���EP�ž�of�iΏ�Y��̐kmF�GQ���z|B"��-��u����[i=r�'�z;TA���=��O��P�;k�����ɑ��P�� 9�Wp�y�O���Zٍ������~b����0����I�cV-���O80Is*�k������L�$B��G���V�����ʢ��v����/�2#��l�)dY�?�q��|�LT�/�� 1huN��$ʽ��My�e�型�{_�E�����kx�4�	�8g�M�t��=/קS@>Ozג�v�%���d�e}�}C��m���n2�c�X���v��8��S�_��<�����w�E�<��c[I�I�$��?9F��z�Ւ�qC�IΥ]�#��j=!� �g��Ea�1z�|嗎᛼�U#ؙ�d�H���ԃ���@��{Uf����ai�3���4��ޗf�#m�K�C(O����Tg,&�ѥ&�E����e����,a�Mv������yl�Y�Ws���P�,YW�_R�e]�[i�]�L�ʯ�U�,���u;�R��'�O�Ҩz �l3���_���&G�n���%EN�t�ƻ�t�����?D���V�w4r�k-t�ub�����RG
Y�C ��y�,R�o�8!GW�2��6��>W�䐖���aΛ#6�������
S��D?:�M�*:��*<���O��ij	�]̤sH0�|�2�wu�g��"�:�6h{X2𐑴���1Rh�us~�ߏyBe�'8�{�����E3I�.K�+GeL|�	��ca��K�|��@!���6������|�pR�A�~����[.�i�A�A��s�W�x,�$�'jtu�L��
���s@������Ӎ8�~QTj��"�P�\�}��p�,�k�痦9=���Z���x�\�%^' ��/��Zo�䲨0�Њ�&����j��z�u.�亓ȥ�:�h^/m�x��̾<�Q�z-}y*��F���Y�*�@����&�tt���g���4*����+��qM��~��ͬcn��g{$�lT�O��=�y���m�Y6���%l�����viG�K���A��7��SMe�;�Zhn��י�]�
�T�x�"�^FK�)�.�2K�=΢MiBl����}�j�'t=�EW�j:���3����1�в�z -�ȪPE��_��H/�E�;���D=��yF�}�%+�ގ���wS˖�L�F�������!���������c�#�]k���ᷠ5���r�H6$�q��(��
�!��8�)�@ ���>�i�+=ho!$D��kEz�{��{��	�6w�G����(��ZU)@�	a�Q��Gs�P9�ϭQ�F��{��,^��i{�.��E�~ "�ȼYc�|�lh%2����hg�f�cڂ��`�[��4��	)p����I?ud���O:ɚ�j�+�6�_�~��9OT�l&F���D�cZӌ-�2?����-��K���,v{�5д�	e������Yaf�?�V��Σ����K>�1dK!��Y쯼���'|�Z�X��_$�����7�DZ��$�v�Pǡr�ߓ�o���#����{[^P��b�\��h�/�7�?O�ymG�}z2��Ɂ[�g���R�>]����>tj_+̷s�+�RW��t��Qp�U�B�?k�W U&�@U�	&�P��ҥ��T�-��\W֜�`~��X�.�ϖ�:�W����x����5�̀���e�
kL����SZj�N���o�*"�/��p�*�),��x��52A;s���ۘ���`��YC.\��<�o�&�	����.���	��}[��M���Ar)������>M����p��=�e%��A�5	Zr���+�G'�c�y�
m��?#)8���w�Cm.���.�m�Ѣ��! S.�_҈�{݋Q��::��)��ϡ%�b��ٮ#��r�U&rv��ش=��P=	F�J戀Cj�'�N�u=�(rg�SUb��(d٪N�"�=�;��*m��=c�V ��2���U�����k^jT:?L5�����?�i�Ңϙ���ć�h FV��imߖ�`@^f����V�L^N b��Ke���b��b�ļ��/�Q���ov�.Um|��kO�h��@��U>�Ͳ÷��j$~�̪��㠚��㺂~�Cp�F����x�����֐m��<��$�t���B
���#�G t&�P��fD�sxX���J��5�\��C�ԓF{�Z����s�d����_����Ma��O���ƙɢ��ul�n�v7D>����aO���Ye��d�I�����ì�s{�p��h�?ˢ~�� �ve��-�q���h)������V��}Ta6=� �ol�;�n*���e�+}o{�J���rC_%
[�/<X���q�r���hyx�z���_{%7�QC�&z��J�@����?��<B�NC<~�e��"TRJ}�7�����Az�A@�Ӏq���ܸCv�20`��3���I�p��!��b��\�i`�>�א���%G�q��F�)g_ؼ�ua����G����������ÿ����%I[DZ�7};�I��=9ߟm�.`�#R�����*�AϚ&`	a�F�:�e�G3R��E8ݳ�q���r��]�w�1o���h��OuO���.�a+I��9�\�A�4u�#�=ꢽT���b����6��\ms�_���;� �i��B�,q�RB�W;Jj��@���f@���B�iv�Wg���BNp���J�-�$���_��Cf�
tJ|�F�P҄����^M1�0���wg�%��zܦ��Z)���f�"���R-�����9�2�`�y���O��s�L��/�_Fh��]
t�'$��R���8�=�`��z�4���r��8��#�D���P{��n�B�|���������k��,���w��[ i�M:��+5G�����K���rE?�$��V��5p*]`Z�A;|������p��P`6�isX����Qe�)�X��3����o�_�2��m������v�P�3 T��;nV) �Z2��g���	��`q�~P�)�CɲL7R��:s�q|���T�Qi�3[������!�wQJ�bO�2o[�O[]ʞQ����Qf�h=ϔY�B�����?�	��$���O6玊�;n�oN+U:�e���V[��hR�n�?`�#�>-Ysj� /��*���S�f�UO~A�ˠ�����4)��gv���2w ,L������ڟ�[C:��|'��'@2-���
fpA�%�����G��'�R��P�s��`��/5���a����#��]2W�
D��U�v��8�_NKO�����yE��5�K9~#�22h�>ԗ=��:��Z��^�$��O�a�W�l�30.����=	a��{�!W-of�E]@p��}F�e��r�K���ܺDIv�A�f��Te�q��|�rޔT�V�ۃ��\rK�U�nP�
�9���h�}vk����@d�;�u�6��a��9�'O �B��O���Rp3-�]|�>}�H�跃קn��{�%ʧ���ҦS��NT���%�Q������Zr��eț�HX������ec/�k}�T�_:�n>��9���u�=��]&��N������f�V~��4k�,3]pA�]��e&ձ�i}��JEp�q|�0�����]�����EH�N������ώ��ǵ�g5�>=�d���x�L�UD�
�_�mW�^-�5y�6f-4�g[�����Q��%�h+���EaAe��6�����&�s��1�7v�ڙgt�O}*��P�'����V"%��������_z7[(������b~�^��|�T�.��;�7�MG�~�����t����E[�3f6/��eМ��K��� ؼb�w�%�Ȏ�ƪ(l�LMi��ܚ�F>�f��bR=�Y�!Z$��j��u�/�zE�hL)w�Y�g@먋�<t���r^���i��?b��g+��a�\S j������e�"pL���\�1��S>��m�)�A�8s��^�vNx�J�!`ژ��������ȴ��Z�K^?��㌍�,_��7'^j�Y-�\-Y�;�F�7�!�q[f��sKl�l��;)h�i�l̅��c<Uȵ6�Ui�I��kh�Pj����p��m�T�x	�;A��)b^.����Uc
�S��F�	Wh��`{W/���g�m������"7��&_<��0TP�d6�R=k��p���o��ħ_{�-����1=!���	5���GX�����)pܳ�ZTR�[�X�s�/N;�N��遥�A�.�y&JT�ld4�vhW��\w0޻�sa�S�Ok��0?UL���lD�����~��Kx��� o�)�l���9S: ����N��"�<ue8�x,�q�%���4������>[�k!����t�~SÕ����=�0S�MtK%6�$'E�q3�d ���v�-�Ո�4hǇ���Z8
��@9��rp�/Gdyy�SU8]�}L��I����.��B�^��{�`Oc�i��Kxk�4P{C�]2Ǹ�RX|��Cwj��dr 1{2{��Yf����T�[%|D,i%��N�$��k�žj�sg�U��D$�տ^;��9�)6	�b�p�����^��w����1���������N��#���>�5�_�O*��=��8���%K!B��l�����$� Ϻ	H�*�۹,�J%���R��z�ҨK�Ƞ��߷r3�*��L؋Ng�xz�8��_�Pp?��B=�5\�lJņ��B'��S�S�	oa~���9�W�{�9���YΝg�a� %�D0��Mp'��P�`4lJǣDa��=|0Rjf�"R�M�R߽+��`�gw��x���g.h�c�BLX�H�@�ދ�E��Wz�
�bCK�~��y(W=�	�Ea.#�=��GE&\���߈�2;_xJ]�|@�m�Pe[�}o5��
���1�0���([1���T�g�<Mo�wMi�4�>��V9B%���c�rA���vB�c�<������ā	-���A�~��F�cP��i�D��)�3@&v�������y��Q�� �,��q=���%������hMk��r}��v�<
�����<5���`� ���ٸ=�(sm TϺ�+�op[M���j��2CL%��Gx��`$
vM}�b;v��
	�y���*0$�.�%VC�5���P��r��߼�X�2�&�`�����&#m�/a��u�H���|���rpn�Ȕ����J�a3�Q�^�!�8��R�c��q�j��q0~�,��Є����m��؞|\�=��^1�����i���iOJ�t�7�v�C�q�}-�c�8�!���'�&�P��a����Zj�
<��T���M���f��ߒ�]����9�ѐs�|SUB���F�9��!��@Z�>÷�����Ӓ�:Tb"z{�6�2�b�$�x\��`����R�K��{7W�&��Tڡ8	bc%�!3�2R����"��z���s;��"���Ay@�E��l��룥�O�ME�w��|?��'��3)	�YZjQ~��r���x+�z��>EJ�}gwe���X�>ɴ�L�J6n�����v��]��@�J�y9�����o����_g�b����������W��@�uM��c8��8a\2gw45�K��`"���%�ַlv�X<wUľ'�#��%������W6/O��2�I��4w MA:V
(n�1:��f~S���?�jl��J�cvsEWI�=�C��q^��x�����0ke�Lz|���O*P����q�f�� =F�fU�zsW��#J�C�����s?������J��U��]�'��{x�����DW�j��#��\�t�CU�!sV����D����6��c�!�����l��6D�9��O�Qj�w���M�B.�������6��VU������������^>�*���Y�Y���_�1s�_��H!�"̩nN�"��\L��G ����x� ��W|���yv5���1U��v�&!T7���(4�&0
˜?��*(X� ^�j���䣭�ʺ�{���k|��=,>��p�. x��	 D3J�-�	���Pu�I���irT�0�˖��:o�<@�>s�,�Ä9<9[t��ϤWo7�jAyX�+Œ�3�\���:�ct����JQlL,���Ľ�����a�H]&}��Z*U~�qW��6����_,� 9uh���,�M��(���P��s��c� R��GW{[g-�ہ3�l,����|������9M���\��
T���9	>j�$��m�s�8���YC*�L"�[���Y�O��-�&��Gs��W�C�C+����)�$Vj�0]��"�1�"��KHS�%���c<���e-��q�>�y��	��/�N���@zMo���K۩y�4�͞��i�W!5�^�\ϲË�H����Н��x��ƺ�/5���O���
��/t1��y-����(�7e����n���g�։�q���CA5Q�Z�jFgjN��9�:�=tƧ4)D�u$&ǝ��F|"��kI[�^�W�O�����Pڤ|M�3TY�"�^�Z��Ye�'��1����}��^S�]N�5��8s�'��
;�μ5;��=��Нϊ�
�rK�z� ��d���%�$>�o��F�ŝ�Ҁɺ�ى���2i��>����;���7\f�Ť/2�Y�3���J���՟&�E掴�W��-x|�Eϋyy��"QB��7�bd��{?/�WNL%���Б�Q�Zbdy;k�%�ў:.u��"�k�ڹ�pwz���A�:���ٛ�N�8��s�p�O��l)��[Oy����y�j�|e�$�)����4v	�f��3�"���}G���8w�7��'Xohmiĭ�$�Qk]|U>B�1�� x���˧-�����]'Z�h�3Hmj��{��=�[����N��?��:-5[��N8�^c�ޏ�/81^,^D�7}���lb+���$���bo����������n�\�qF��S,�e����6|�W	Y�i)��9ޑs5����T����2|���L�w���z�&bo�P��6����Q���i���E�$��Y�c�-�o�_?R\�.�4Rz�1�IP�NLU{ބ\�|b:�'�H��_�nWM��yt��9fy�� ��h䏥���%�֛�z�ŵb��;�vN}e�|�],p��K7���JuKM�VI޼�{<-{$='�����xS'�
F�gvA�I��E>ѫ�t?��\���|�>b�ntS�lFFĕ�ǹ�7�j�hpi�q���b�>{-��
UA	L��:6��:$��8DC��C�Gt��jL��h_����a�n߶{G�JΧW.�z�ֵ�˱}H�Y�q��L�����M�M��W��D�--	.z4{�V�;9׊����U�������F�� 8cZ^>�I��J}��z�Y1��z�Q�-�Q�`z���&���这pl�f��zJ�00]�!86ߟM٬ǉ���Ϛ`�_p[E�v0��ׅ��E����"�6P���2�h|���G��.}�����t�p4�e������YU�DK�:^�W�<a�}g �y��n>5�g���s*����I�*�������-qFn���ܫ��Mb�;���y�4@@Ǟ�0�ay��d֯�/��_<rT�Xu�q�jɋ����MpvJO5���s�Al���� �}�BTǝ3{����L����=P��˝�����
�,Z������Rj�����5BC�"�T���s���7�u���	K-�i�C#���u*�Ƌ�?�"�zQ���2ί��̪������yV�ͳZ���{����W������o�(��u��-<��U����/����zV]���U)�u�v�B�B���,b(R˴?���d�v�i��ɾ��z[���*h����ŭ�l�ȵ6�~�qQr&ȮWz�e���o�_XԮ��"���3�t��y8�aQ��斁�OoRU������*U�ؗ��0�z<��@��~���W�]����>s\�E���TV�s��e�|b�<�|גW���y}ZӒ�pS��v�4'�ݠgMx���y��au	��hhM�	���+����Zq�G
��/(ϙ�v����֢�|<d�)�\�T�z�w���g���#\L����N�6�D�L��y�W-�f��Z)���D�2X;�|���{Y�[� ȕ�9,���J��EO��z�*h�.� �y�_��(�Z����F��o�v���O0j��i�|m��z��x�m�q��܉�M�zl��U?HfwW�蓀5���c�Q��Ҝ箝m��z�Ǽ�Y��6Sp�>��}���HI�Ti�
r­��������_�;�e�WZYa6!Fy9���#\�{Y1�17����g���Mg�7�E�/(�#77M�&d�c��	O������z��x��(ޱ&��
-!{�W���$Ĵ�ƚ��'%RR(����){��k)������L｟{����?��O��6��Y��~�s�������5�W��z��ѓ6�� -�a�ܔ����{���(KS��b�Fl�z�mrJ�q{M%L�-����/���-�0�j��5M2�8�S���%�n][dLff߿u{.��YAn�I�?�6ؚ0����`iٴ�]��b,z�8�
Y���k�i�h��5��X�� �Ajf�`�o�.ٹ1�XF�m��a���#���l�+]|o���
	%�4�l�z�66�;�v�P=�o%s��j+a�W^/%�%Шs�>k�W��? Z��Ģw~~�:`�{��3�;ߊb	�[��X%TS�~A���x�R����q(�h�ŋ����&������� W��{.�|�[`��3�yL�2�}��}ѹ#&�<�t5C��V�Bؓ�$��E�~UT�� o&�CFt2�s�3�B}Sev�`�TY�ռ	6�����U��q�S����;��ױ-���sѬ8ׄ>�>��Tr�(im渗vˍ�L��/�����9�����u�� � *_�*��"�m��Ӧ#8KO"�8�tKW>T��R���`�J��H�X6��_���(����)jAS�ܵ��l���*(��HZ�]Q�L��Si��{�`P���wD�o� �P�.C(2����^�VM��>�.}Q��rgoüp�:�b���,�(�'�LĽ��/��W��t�"1f7sp�V0r�;I��q����kl�HaUT�^3g�6b{zk��f�A�7�����h��w8�[đ���V�O8�u���5Kl�f�u�^�f"O�d]���]WԔEض�?���T�Bw�Ҽ4Ǫ��V�_��R�.#�d��K
Ӟ���6o�g�����?�8o_4K-c�R�Ic����(���Z����/�yc�7tH���ep�T}�a�����P�c�xPq���*~J���R_u�Q����9����]����'O2��q;`�~��k�U��B#��I�����"3����	\�=F�)NW�|)Q�\ާ �ewF  5/c�V\��C��o9�,N]����zZ�͋���|&V\��k�G[+�H<�]��KuF����F^���$� HGé�X�vv�'Ϩ|H�.��z"�@�>���+2ct[�dz MP��Y�Jf�y�)H-(�o8�������nQ��Ɩ���t㪔+B��k<O?��ߋwHj����"�Vن�����(!���)Q�~:~Rin�vK��)6���F{�8S��cU6EfL
���@��^��m
�L��5�;_R��&7/{-�T���η�eq��cE)c�Z���
�[�,=�����4j5D��e��c�Iu|�ǒ��[~��9ҺB���������hA�v?U`tC]<|j�����^Y��Y���c}����h�o����dV�]k�/��ezX�S�P�0��S�G7�s,����� � C��AP$�����������,%y����g�G�dl�6Վ��S#�xf�ç	�n$��D[Z�7�\�S�IPTkų�V��<|��
�0;9��F��е��!��:Cd��F�A|�������t�-�Mi����p�t���}�a�A�>�*	���[�} ���"r� �{:Pl�C��2�
Y�φW���H]�񚠠�
�� ��+�:%����Z��f~�̦Oפwu�osDniN!<[��	�1>�� `,��~��5u������'�.�ތ[�w�{����S�J �VF��^�=/]���/asw��㚰ar��y�O.o�E�Q�Yq�6�^�%�s�A(�M=�cRzU{���p���f�����+�Ԯ�l?��#��Qq0��,�:l�@ٖ7����T1)�:ٯD����\�*D�ͱ-�c�OA�&�F�ډ5�&1�+���3Nsy�P�����:m��nM�$�E�oV���M�vF�}��Ø���;yB�X"�,����_��?�U��dϯ��E�����GO����ޫ͎�"�O�������0#�G���G�#gӞR��w>�&���Z��Z���-��4z��)�Y�4�������7��6�`�����&�_X���Dk?"m.:�u���vZ-��U�zq�ܨW:b��<��u.f��]բ�[��¾@�(}^��8%��m"�-��Я�B��ⱹ7�B�~]qe^�<�o�HVk��mV�qF�}��?�.�����x����L�>��!���?7�T�﫥���<�-4��b}y�U���['�5�Oڢ񘈕�E��ʇV�y�ۿ�m3+3�u�m������z�ˤ�Uc���ؿ(o��������zdf��(aoJ�`&���*|	&<~R�ռ� ����x���i�@lfv���GǑ
�JAn_���3H[�DmS*����*{�b�VZ)���"�X����-bvo���P�"2�z�E���v;�v��Hx�}��`�.�6���q��Ÿ-�%�Aj3Qj(^��!U9�}ļ��S}wer���m��Q��#>��
�Zo�Xk%��Mx����/K��6�<m}җ�=��6qDm)'�@�=�!{�!�$�xA�j����,d��ˢ��T1E&���#ȽV\��Òi���x�{����\
���M�� �a=�5QA.�/�sl}��'�V3�C��M��'pδ��#�0kg��ռ����«���f����"��t��-g�����R#"Qdn�lxN��
�B7�~�u�	��}C�s�$�ܢ4�����>Rֻ�w�������aWO�+R����y�w��f���<L/mN�rz��j�d2�3����.�����r����n7˯�b�(���iGΥ��
��%��E�i'^�n�8!q�h��G������~U���3M,�UJhm~�������?��q?;.�eA�������*��BGX���O]v{�Q���U ƈ 8C8F����H׬���t��0��r���\���;���C]�{�(_���._`�),)s|���S���ě1y�?=Gg(e�=9zD{<��+�c߲����MM^�iQ:�b�"ڠ#�h#���ۑϋJ5���i���縵*�m^��1o�������6���h��E}J;�ac���`u�����"�� 6n?��P2�|�A�fn�-K�j�Ƙ�մ�Xm��d:'v6<���1�N�1��Q\��M����Q����Z�����?g�3������y���R���]YZŀ��I��>x�o��'ɉL��T#"��|o��攻m�xV���xx_�fV���L�s�Ӟ"i=�z��ZԿ�B������}Y�$���C�F/�{���&��K��y������%�����n(M�-s���[Ne�K�����֑�E���w�ݝo���"���c!S�2R�\��sL��Й%
�$X����,�;��6�h��yPb;�)��b�1���V�P����7�	��S�����
t��$v�c�T�������x�
t��JLT�g��L�z�il��H�;��{��|�݋
�|fIݢr�D�sh�'��V�MY�E�S�	�c�H�˟���-�y���Ηy�{*�!ޡ�z8��{|�8�8��/(�Թuڟi
��s#�=��Hv���#�2��(~�;����@�xql�L��G.A�p�H깝��܋������W��r0T�o��-� L��qђ��[������s""Z���0��j��#�I�W�b	>e	q���Ǳo�3u������wd���x���`0��3��9qy���u���ˢtإ��Tܴ��d[���*���D�ǽ��숾{��*����x���ǩ"����f��'�nT��!��3�&�l7���__�O�w�r[��)}?~��YM���Su"��e��L�) l�Tn�
oI��uG�ط�P|�@��nOS�Qk��>A!��c7撴e�\V�w-`�*`��x���(�gp�7�9��:���%�3#"�)Q���l��^��Z��1`���Y0�amPDL]�L(b���;���2�~��,�*��i��m�#�"��-�j�[�S TO�b�oo�U/����3��W�_�8K�;NM�OS����(B�G���{"��)�	q=��x5���#�CK��F��G���U�~��<%�;Оo	yQ�*E䣪�Qc��g�%�`�7�o��nxJ������2��z-���i�B�=b�׾�ѕP����m��0�3j�-R�Gc��N���(4�0�����.nno�W ��q3���à}1@
��:*{Pb������j�{��G�ʒ�B�ۙz��6^��!>%_�J¾D���SDJ����������l |�a���o�}6���)�X�Y?oa�1`9:;��*��)�"e��F2�jW��:�^����V#�_� � �i���Yr�q�Ӓ�{~�=}f��k'WҮ���l��$�)�F��}�6�j?\���9]�O�� ��]����Xq��++�-���]��,�b�z��yp�"�=�:L&(KX۞J/hqW�L3�!re�=�m�0{���~^W��Զ�YW�_A�L��L��{�9��`�a�T��ǀ��7�0���Y/�j�3��(O��IV����3V�HȿҀ�w+ܰPtf�w�5Aq�L���{��k]:�0��w����xp���N�?;l��P�v8jԲ%�|ȶ;��$�n(�V��%���e`�v������fi�Y�	X4f)��?`>X��թ6O*��z��ȁ�_�9�@m% �v��'*����_\X1��udM˃l�E)v����;�>���45~��	�,��ҍ	ҺW����4��bQ&W�L?K�MA�.��L�1:my&@�zǾ�ycp��ƨ5��&i}�;j�P���4?���'�r�'�Y����`�Ӕ���4����`?# R�w�ú0����6'�K�_��x�� s�a�!��W�J�;�(�k����%��1��k]8���.�%���S�^�&�N�X�Nj-�w缁I�O��#Cz����
ӎ�mu �?|��~��!9Ѐk�jN#��|�ӫg=u��3�v�������S�;��{	p�p�0(�x�ۅ���������kQu�x�,혊����}�u��X&��ӊ�a`�8;HN�Ql�/���6�#�*O_����"��j�g����ʺ������6�8�70M�L%�&wؔ�
�n*�)�����p���$׬'j�Z#G�g�9��bՖ�����8����,��7Q��7|����Fd�r=��D}�Z�Ls�L2�IuO�ޏ>��(����^���79��#�ejca�xI`D�c�kbRޫ��F�YL�Ye�-!0�q՛>2n0w<�����U9`��f���N~?�}��R:�%k����Xo#ו���YI�&�}�l��{�En��ʍ>�e.:�ܻ���
R�v�d߀B,J��ǯ��
��zĺ!� '*�ʖ��6e7�(b��)
�;�����;��}�L�ٚq:������O�R�_?�Uh��'&�>�([����k�&���s�_��2g`�.����cK�Z�0�U.Չ/q�3�#��	]��h�H��wJ��t�ʒ,�g�Ĝ�$���6���#3,��2'5��;��L�;YGt����sĤr��g�Y��#��i!2UG�:�Qb"N�LC�W�����Ԫ�g�b��}�{Ww�n�e�'�m��^�:5���}K��c�F�����`�}����I+I2ی$�h��E��%g��>G��1s��1/2��߂Q&'��f��H��� �З�f"�DI3l"&ó)i���'p�����[�a�>��V��z�-��f�y���f���#�)i�A����2D�޹�?�Z���z��[���xt�]Y4�W��ךcx��ղ��_Ѡ��%�od����ͽ L-������_�Ӄw��a@���DG�e���j�uu7<�o��Rph��iKR��������F����*4&��2~q��ζ��T�	���R>gw���C���S�7����0ζ��}[����B�Y���xW[��\�V��/2����!����h�sI�)��Xo�9)#W}g��z�_����/����hy� aߛL�IMYkX�Z3a�����u�8���!��0���+���Ȝc3*gԯi�	����tG:����<�`6��us�M:�X��z��Yؤ�����<"���O�L�;ͿL
5����!bV�So	�0��ℇx�jV���[�������i���5X�N�a��V��U��gd?��B�66qߧ���]��;�.��˷z�ScpH�SŞ2":�<h:R�SwBf�1?����mwxx�*��87�(����'����o*tTC�G�WD�,d�V>��<��o�F�h�i��h���(ݯA�Ŋ��;�K��j�|!y=<�F���1R�e�u��߅�d�]{ER�R�GN]�^G��x9�#qNX^�q�?*��L?����lI�f���wW+���݂UgB������;{�c�������z%D3�������k&�Z�,
�˻�"B�Y)���d# G�j�.�*�laoA�����^R�B��$�je�w"@D��Nm�bYpN �X>�E�׊W���%y���=[.N���ϊwl�\��Q��5���
*��,�_���a�U{,��>���tU��~��w�˟�,��Z�S�ϫ��xZ�Z��{ۀ����|�g��7��Q�~ź�uH����$s_z�B�F��f�pv�˙���e�a4hO�,��RI�]D@�$+��*�|��+�aG8Gk��RÃ��ϘxO]v�֑����:�������Y��fk�{4+����j����;R�Ah?X�ϭVu��Èpy�݄��ȯpI�b+q	���:��s���z�tHo��j�Ò��G��,?%��ˠŅұ��ԕ��V��>iz���T�tk�=-&���e���+r{�]�le� ���v��0�g�gY-qd���w�c*�Ӥ��� Kz_�@@6�:����s��>&��Ot�ʰ�x9�"h�Z� Ȑڎ�Q����f�Z�I����|d��#�,�J ��F*�lƿ/��~!��4FtA ~��5�e��+��qӴ��YT*�!c�qvT��~Za���k��yP�QjQd?P� �j_@����`��.x��e�����{�4�nj�;� iz=+)��l�ɮn�
�@}�[#d'ҏꏴ�4'*x��2\1s+#�����osn]Ce5\^B��`αi���c�Mm�8����k��6�#%L�^{��X��'���~��EhGo�/�}\��׀A�j\3�N��f6/5�i�ŋ��� w6
�1d�ƽ��D�f�v�`4C��ơ��7}��=��J��Jb�
�΄�(��O���_\�;/3O��Y0�U�c��S��5)�1�ޛumS�nz
ȶa��X�M�B`wm���Rm'�i�gj�|��l�F����m1eiJ>ص��w͂�7I��9�4�G��TJ�9��m-_L��*�P>��f���6�캂�P�C#:)���T�|��1,�|�D~6qoÔ��[��3
�Y�1e���{Pf�]x��Z�bcew���>&���ذ0��y.5Mi[���+��v�1��!z!�W��o��]����㬄
�L���	���(�7�{�=�
�
�n�+�p�p5���+Q��r�9&��t����+�1�l�O���J3��.�_������a��^����`�\r�};ٖ;c����=��o���q���=����G�Xg�u ��n�ծK2E�/����O'��uֺ��<rNN�T�W<x0\d��A�ί���ޔ���2�$}�&������Mu$nO�m��4CiR�/��.�[�\����KkS~7x�[�u�m�~���!��$���`��d#���n��ۘ�B�g��pKЊ��鳾��O���w�g�ú��"s�~N�D߹x����2�����T���R�;o�p�Z{s���y��cf��>��q���$)l&;���vf�i>G���<5�`w��j��T7��H.���ڙ�����\
�\�@�/,�kG��H�bl�!e����M����o��23)!��K���S0IH�e�0q��!��+�P�����_�{�02*�Ѯ�8��rM55��x'�̾�9�2��$
RZ	pD���E�ckW�éF��9(��_rJ��J$�im[���ا�v��}���\�K���R�G� ��IJ�&�j������#Ȣ'i�LQ��62D�æ�Wƭ���4�\��P�N�'�$��I�K����0ĭ�թ���ZΐQ�Mf���H�~ݺ��:0 ?�z�Yf��ŉ�F�E�����Wٌ$zO~�E`����{�KI�����<�c�Q�\�]� ǽ�0K�_t)�}��k�[��܍Н+7LS��M�2*H���~��.�$.W��_9z!l_\w���.o�^�uN`
�nup�ű��~��7���\�S�p��=�ltd�Q,_����f�3z֋���#�d�Nq�o��	�L�ې e�^��%��=��ȇ���
��[Ik+��V�dbC��o� �t��״6�Skbkc�<�K��_�Oϩp=��6�~�"�r�Q�H4�j7�`$Ᾰ�s�����[�V#�E���9��Us�¯����0�������;@�>qJY��Č��E#]�f��o��'�v�Zl���w��6플p�&�z���q���X������߭퀃� ���`1�>��/�Ȣi����{<���w�'�U4\l�:C�}��w��|B�:���ru�Oxv?so������Xl�K���,���Yk#f]�0U��WBi{첼�J����Qs���UQ0��P��8�lk�����Is�"�Vy�V8}Ʒ��P1)���m/�W��QP˩;�M5O��w莂��ak�c�`����ѻw��X�/�o�O�%�۶;��g��/��������ظ���a}z5GCE�9����? ������&�b��RHu�����Q�A��� Er�?��	��~^�l(^|4W��̐u��z>��Pɴ2�柂���R�|K�}�m*Dd�V��Cl�&���ǈ�)���Q�д�9��X�"z�����\��w<w�����bZ��w6(鼈@`kb����v�Q��D�p/O�w"Ε.O4���(��̸��^=dD�0�lWhR��o����5�`U��4���I��eM���_rN`���,G���7������"˖
���X~m;�2f�1�<����$��o�&�wg����¤v�/��ќ�H���\����\e�4��:h
���w�S��-ս�F�E��x�s�2�J�h����ճ�nӺ���~T������idh���A�><�T����oOQ�X��9t�am��O����.�F�w>%A�޶�!^�IYg�3����2l,Ql���Y�u�,�#�,�K�~���%���u���\7�>�s�VO+n�����Z�xY�41���7 t��Ң=�绽blbדoڷZF_�88��1j⥮�9�¾�[��&*�5q��Z�l�S}vv$I}'�5�D(��$N!Ȍc催^���+.�f�Q��-�����ߎ�x�� u��Z��3SCɉ�9D�
nu�`����W0�m,��B�H��K������8�Kh]�Z�Ƭ���@R]�,0S����zn��v�D�4t"<䖱�>eZ�OP�:#����mV��~�-���}��}&�݋���(���ÀԚ�Ʊ-�Ftv�<Kóؕ���|9RP��r:-��=Pd��9���Z��g�X��kn��FRX�Ŀ��~a��N}���o,�I����	���uŉ@�~ѭ�������
m"�۳�Ӻ��o)�����?��g�ģgv���#��B��g��V�j��ͿP��⦙��<��-p�e)Q��C�t���oDIsω �	�8�-��?kCDEE[+f�������}%����-�?m�ciX��іyW��s��������� W.����!&��)�� L��PQ�EH�;���|o��U��x�'����c[Q�X�L���%<�~4��[��, �����;O\�=�*t�յG�(�~���=+���JeoFG�}�0�Ɔ-�+o�^!"��� �#��~�S<r��
�za	[�+a�0U_2�G�3��3��s��ހ��T���y*D�c04� *�!"E���+-�����Bd����/\��`)q$��]nFM<��k�!��0Z5���fp�aP���q�ѓ6��.�7y|7(�t����
�E07�6����׎�C8�����ҩ$��c.�,�;�'S�X3>1]�����*sN����5����3�lj"P��i�V�[3��!M�V��Z����JquM��9�̣��V�>3�Dd����&7��9@�ܲ�����:z��ƍ1˛�EH�2A���7`m�lw{5y�@�/�wɥ�Ϗ�|%R�6�*�&�Ow|��j&�Һ}�)�КAɖ����ąC,T���#��n����7���`K�4�����P����b�Ur�w��??���h����82�/�4=��M�}�N�:¹ޚ��P�na�S��xckw)��O��O�oa:~/�?0��!�\��SX�rm��Z�@�s�
yV�]��z>��p ��>�L���T��	o�H�+��塴��D�ã�}uq<|�p� TN��p��G�q�][�?'�K7����@����^�p��o��f�o���� 8���QP�����4���B;r�N�uv���'�_��G.�R�֨��$������zW�.+�.�w]3�&֜J�O�ǯb& ?V�%'�Sj����1?fL>�T�F�fKT��J�C3���٘_^/{�-v~	��D.ǵ���\2w~�n��ss���K1����Hb�E��
_����@�z�:T�B��6c0�-�!cjNhp���x�#)0���gm�
Ĉ��wf��%�:īw�l�Ń��]�t����#F���U��YM�ϼ�F�~i���1`����0���X[��6�H��^�w�l�SQ����Q��-��El����<�G�2*� 5��T�b��i����o��rt�@;9$�������&�x��8򑡂����s}�|���ޝ�S�R�
�0��K|�����*7v�����>���rؙ�-aD��nY��+�.��\7�8�Mji&ȟ�4�Ӫ�c\�y;:ŏ[��-\�'�n����3F�9C`�8y�*��������#׫�H`)F�y�W�������;nYBx�_6ɸ�H��"���o��+�]�yJ�����
;��te'���3]�R���Q4������4�*����@1��r��N$�/�+Vs��<u��f�S���V��������2��r�+'�Ψ�t����P� \�ly C);�hT���
�/m{r-��/"����5~B��$�MR:̹�a�#�}���qAmi��� �|���;�y�5b�`2I�ﵩ��S'Br{�B6p�<�W����]i�^�ݚ��P�`d`@�q��E��lSaBi�)N�,�"���S$��oj�+K��o��k�\��6��_~���z��Emo�:ٴr��5�>Fk��:n�ww(�?�����'�����>�"��u��kޢ��k���i�K���.�g<A���
�1W��[��_� �%��Y�h���"O��Q
��gn��?� Ydq���b��tE���L'Ypnu?j�c��%�>s��Ct���l�Ja���*l��Hh� ��4���C�|/��Q���T˛��q<"V�tegw�͏�	��Pޱ����j����0�2���2#�]5(_[P��U����Q^�y��hq��l_a�̣"��aW���3�0�0)��$�$ �Io��تgq�؄k�R��_�20|�IͶ�ڪw�}~�,��m�)��i��d�ei8�]�q��am�C�P���,�ꛦ�� P���gG�.g���񥁇�ƛG �mi�}�G��=��V�� v4�< C��Ra�%+g�����|#�߭o��
rv_�;uû���ض2�
���(x_��Q�R�l��;
��v6�:�o��e��A����haX��]_�;{��Y�_(y��f&�/�@�����ac[{��̳�v�Sr���/��I��������`�y��^�g$�JY}�t�������0:-k�{a���B��"����-1���^+��"�?��x����O�ɐ�z��{��ɰ��%�!�u1`�[��e��5�{���:�g��˰�@��O�9��+w/�����z\��8��<Tt�| D���JD^Ӳ�b��F���];����C�T=;�PK(��h\�	C�y�"l���s"K������C	?���O��s_�y \�`_��Mo�T��M 0O̷�TXj
e>�-K�q�j���Qr?��V oN�j��m.�D�2��g����Т�̉������~��yi\mn��xo�E���^���%�V#��^��!_�}� PUy�'i&��3*�m������Q�aa>��\ǱgW���6`���:r;Y�����'��߄��PD��kW�5�+܋�	�wK�?I��=[?1���Q
�A:�w8`xG���6�!����l�vѹ��l�h��8W��E�;!�5�˿n���ص��,�lf�Ġpo�����&P�1���J;�8%������5�>��zV8@�ݔ4&���� v�˺�&
.J�%
{��w
YW̟1�?�lBn9|�:T;c��B�;�0�h���B�� �8Y[h�G0s��t�v�$�{&	��g��� ͇taN�nߒ|Ȳ�|�c���(�+&i�$2�������_��
��6���1X�������yF��gGOq����o[}�Ns��/�_K�ev�wĴ��������һ/��o���������x8D��=+IΜ|�kos�3cZ��ڻ
;�V�x_���*�%�܏0V!������aS��67�̋X�z)u�&�^u���Q���A:ҝ�s?f��aS��O�BI<�␇{[,��9�3���w�΅�#Ͼu͎�J���L�[��vr�ہ�6�@�C��:t��{�17s��?�㼚:jI?YI�8��;�kk��ﰞIxOn�Ki��օ���џYi�L��3o�|uH��i�����RǑ{�a��w�`?*Y��79H�D����|s�w�f�ۛ��WA�$W���o��n�@�=¶��V��N���e��t}�
h� �����|'dpA'I��ə�7�.k�x3��F7�*r��k h7F$@�U�^��~@Y�=��*�`�&��ڢ\�Yr}lS��mX�Y�.�|��D���k�vf�]��9�FJ�`�E��/�Ӕ�6�t���&�}�|ȡ3�c�!6J�q�`�GP%7�_���a2\���k��X�%堮JqD����R��
�V fM]`l��H���[��A�x�0�
M0�ƀ!A3�:�5_�6̤��Bg�9���b;pϖ�/O<���E=��pI��2���N�)q�[���>��^�Vz����&l�H�~��9 ��B��꿻|#����s��<eo���t{������w�9����g�X���G	>�Ϗ��A���hf�Q���F�J� �þR"ziO�s��M�#7�_�,s��	��ձܙ��07V]ݓg��bV{�� |��(I�'��0���Mӹ�(�Nj��<޿�K��{��4�v�YAj�`�b�Ėh�[{uhT��RG`�1,`��3&�F��5���+`��I�N@��.-7�9K~�2R��_I�*Q�K��I��e~i�b[�}ҜǿcOD�K��O�O�����?F��	Wo[���
� nQ�(X
����q3-qmM�;kݟ�.��w�KS�˧�p���
��~����W)*��$����tTVl��r<���<0_�T��b�����W�}yB���zE�@Ԭ��iTboܲ�b9���K|&�m?=9[��ϻ��<s��=��-u�kW�?�PK   ���XL�I�� 2� /   images/ecade926-82ba-453c-8c81-d3caca9f3c08.png�eTTm�GD	����s �nPja����.�E��s����x�g��ί���Ͼ�k?'LUY�#*1*  �(/'� �� ާ#����l��B�.� �{�{�$���  //������մ���iZ{���"1B"��X6y��z�F*)!�d	B��`�/�g �7����1�y�SЪ�8�o�[���	��HG��fgg�f�f�V0����<r�P��r([���Z�W(ku��@o��i�e���*i�/e�j455^\����]|}��UT"n�a��ww��K�����~Ӎ��9��qDb�"V/F՟Ȫ��k�:���Ǘ�ǖ��d�W�@��;�=R��p�_0~��E�ֹ��f�
ucX���'f�l+��.��-"!�)L�bte{Jm�/��G���'��S�mO.}�I���^��R;��Ice��ʓ+��L0����A��������W)fu���x�_��� �GEذ�)9���tV��`
CF�{�y(��3��^�0���lMףz�yW/��[��t9Z�����e�vD.0ˤ4!��%�CM�Kv�%��~Z�B�NP�`NuU����	˪����z48*6P�+Ư�m=s�����rI���J��^�/��: oC��Tq[�ʸ~��4�}�|9 sS]2V�,6��*�N����7/�p���dcECv�b�%���`��VѪľ6�ҡe����"��v8lY�L�A�D���&|�Z/12O�92>{�Z��t�M
��-sq2n�x2�09��0O��h��@�:��"���?cU:y�w8�4�c,v���_6�*؉�������F�:�k�+�A��I�
v�YG�Y�Z�R��փ�+�FM����T����qy��/�%�~�t��#Fix�e=����^,���C�3�#� �s���}!O�!�>�W?j�f����A�Q�	1}��2�� ��ϟp,��O�d2�$������HV�7()����G11Lݻ����Ӝ��UC 	5���`���F���sq^u��pD��[!����M�=H_��m ��p"uD�6����z���Q��9�U���d�6���us��(���I���$�IKU3������rKt����B��)j��@�)�{�do�8[:!T��SY������]��b�>�c~�$*qE642.gB��R%Ww'� 6�n9ZP���Ϩ�%3l���-�R2Q~�M���ڿ���R���er�*�yF�Y�s�9l�s����
��Q��{�ԣ��n�$¨�#M��	�&��t��C&]�#�c(bf�C0���b��"���J���f�<ƾ��|�7�4��n�y(3R���]f��2���!��5���L���Ͻ+�W�]���5_�� ��~+��&^��F���`�>��c7�J��h�`�־�����V#����0B��ݘ{�䦐tY3k�޿T�$am(?8H`�a旬����Q��c�����rؗ��R����mZT��G�A�4]UuͻO.3�il�	��c�NηT.�T�v��Fs+@�*��j*����y	��҈c�z<����g��e���M�)˂���dw��L.��^��$^oh�����-( �.ޏj~/F�;~9��	1�<,g[����x���uRk���د~�8t��b�b��X��hfѱ�\�sbb�+I�����Ye:˖x�SH� ۻDr�G�0����������_As����e����%��jMg1yK�w����Ces����M��D!n�vTR�e~ķ�?��B�T�o�~�`��0��X�2�'K焕DqT6��$�k|��~���j������<�D��*�\l7V��[M���m�ɻٖ~�(_5���G�;'�s�������AZaFW���Ej6���%���g����N҅_���7��*++����	~{8[�sx���8�Vc��#LϾ��5T�P����R���16:Fӳ乛�=;Vn���6j(�
���g��l�T\�Q�ܱ>y�c�OCL�R{q�Ҟmy�O��v-)�~�~�h^4�f(z۴7j�Z#�<pŌ�Z��K�Q5����G͌^K*�/xpk�)>��9�Iҷ4\e-c�B]��n$!�}U���h!���2����_��!���M������;6H�*.xq�̀2 F���F�G�	�L�� �ٽ��l�kM��޽��qѭ��9W7���h�y�T<5�Yr���N��p��ɝ�M�9�K�0�?g��P�)6�H���M8>s~�Q]�s�Q��}����*�6��z����W�D��Q3Α��Ŝ{0HD�0f;rRIY>����S'6h�w���* uy./�E���g,>�7ƎV ݙ���B-��d�E���ifU�֑��$�ƲJ0v�v?�r��i6��k�F�9�y�b�a��c���?����]�9:i�o&Y�K��{�����7�)���3
i+��t�~
ȿq��'�-$s�"��@qT<�L� ���ۿN~m�]ɈLCD���������&�Z�m?�,�AL�����^y��D11�;J�o��[m����Xi� W{�m�ZAbi��};<��`��]�PV�fm�Oq���������N�7�� 22����ItH�<� JM����r?Z[�PP�0ҞR��tT��97�UdbP$8��X5�V��\��vM�S�ȇT�d��L*�i�,�}���e������ٴ�~ ���!�N�b���4�
��
T�J2/���MV)����L`������7xqC_,��7{���pu7栨̔�N!�>�aE;"�t��pU��x�~w?��ճ�B?���Z��R$�hH�,�9�c�+�>��j-�5�Ud�v��UW����W��k��:���-�^�,�1�r��"�������p���ָ%�e�r0x��1Ʉ2�� I~��ȥ��,��4aj��%�(���j4k�V4Λ��+G�kPz�7�m��A'0ɕ����M�pr�m�ӟ ��LL�V�I)�2��9��g�&�@hFp��9^9�W}F���Dfip�liq}+|7�\ļz�$�ܱsqI����u@�	�;Pi��阽�2�p�w�O3�9l�>����3�sm������bV�	�כ'���[��u�ݑ�Ka�Y*;���S���qa�s�C�\�E��?#��g�b��T�-�cYS��e�QlY3B�-�°��O[�1�����C�����ة����x,�C#�m���̤q�%���!��&9 ��.��Z[�Ӳ�}̻%�&��2�A
a5��_B-O�b�%Q�"j>���\�I۽��;|+;_��Ɣ�$]|3�b��>׳:��[�X��녑�hȜ�����Q����x��&�Qv���u
����G31p�
k\̏����ka�ǫ��X��+��іx����ԕ�ϱ�pB�Iƙ�F���[?j5Y��$����B�(����e�О&X|��N�����V!��M�@�Dg�Zav�V'���S�˓o�D���x�&e�a
^	o��~��kF��$�bC����k��d":U'�2K��t�xX苲Ϥ��YDv���S(/i��=���G_�9e��~��(��=����B�����'W�T��Ԥ��L�;�*��-���\&��B�@�ԇ�~�*�n�ђ�+���hB|	�b��.z�`~�� sy��=U ՠC�H0k8&D�2>zQ�m"�=�ջ������e��*.>�eޓ�f:a���M��;Q���"8'��$�nfW�߯�:�l��>�n?��%�j�s&^�-�_�SHvZ�x�9��udzj�,��+��o�vX�^H�� _B�b4�e�x��v(������36�F�����(!%]fƱ
S���=���Z�`���(u����w�06Vw=�?U?־���^���0q`��NȑM�*�̊w���~��w3�L*�=M��Q��U�����G���:��NE�����7��A�
CC_�D�
B��2h[I�Q���F�Z	�s�����tq2����󢘼ƥ���R�-@Xfψs�s�׫�p��M	H�Z'1��Oc�|�q !U�#��5���{O�����ٲ9�(�Yy�7 �/IK����B�m^��4�C����k��P��9u���ۼ������k��,_��糿o��|/�ԺY��Uf�F�!Y������������5� R�!�A@s��4�]ӼXAx(x��7П	8�R7vlCr�>��M�p�ə�4�ݜ[L��!�y<ue��	�=9�μD�qĹ<D$��OS���a�.�J�������H���t�TJ�wA�$�;�o�|(����9F���$�N��y�(|����a�<�:��f�|�:M[޺�T�⏕rY�<�V�z}�MQ�_�4+`*�����0�)��I�=�)���Z�=���2_���旰|дr
iy����-������FGG��4��Xe�":	e�X����a���Q�܆���	]o��Go�����u�I������IF�G�4WF�Z�a/��p6?�7���Ӛ�o)�Hҹ�^Bm�#|��Lc�~�@�տ8�!�erf)>�y��Z�;�B��h�p��7Y����q+�Jrrv,{YF��<ON)� �߾=�*N�ԣ�?>����>Ɣ����ӛ��i��n\<��T�wi���r.��;�����)�=R�8�&�W��SB����s���ᑭ�����������2D;�jE}|�3��zE¢Z.�P�������.%�4K7��`er.\I�~\D��m-���Z숣n�᠕��T[�O�=���ãdje�_�d�~��ȭ��Rט���F�6��D|�J����S0�vH�L���;[L=H�������D}�����2���c�c��WJO����P
�:�/y�þ�Z���'g��;��Z�u�PQݥm"�S.�qD<�Jɞ�d��9��"��M��nNc)_w0�3'�B�����M]Γ��x��C�K:C:�$=M=	�܁F�~�~&���j���������tG���ZB:,�W��W�ؔ����[>5ظMWn�E�M��l������,��rf����&��C��3������zk���VZ�ӓ��|�����}%�%�g1���<k�s��a��U'����<_g����q�U.��r����U�&7��Z����9�']��'�~JO�OJ�W�%+`U��WRg)StB�D͐�"'Q{����ʻXs��{�uf0���^��~\/�'��x��rx��Y]���昊�g1���S��f�	\΢<��֙NZ|�q�A��ih��b�3M2���&bI��+�̛���@�lG`�3[��6��핈~���l-�=��NG���s���H�;,�� Uԓ5Hb�t�q�=<��	�,^��!l� ��	W�K��ʦOt!�9�����VǙ�cm:>���e�M����l���M-�4�ȋ�W�;�j��sT��s�f�p�OXVJ�yQ�A���: ��w�9]���ܨ
	��4a@�ban�Ն���|}�6m �`^�+E��swх��ߘ $���f��u0�i���1�`��~0w�����(~�l��\�*�!�2��D�h?g!$�� #(q�S���ݩ��6�ݫ�ZB�I:)�@2~���@[/R0Y ������\ׇ�n�����K�̴��Mp}�����0jͽiJCz��{<�m3����O�R�����,�G��YKiC�{;8�Q^��x>d��t����y9�k'%zc�F}9��%�d(ʉf�� �4\�"Ѭ1e�TL�u��D6ķ��3"26$�%��)~	i�]ɷˌa��Ł���j�~�#c��d�ꈋ�����J �la��N5-��o{�u�3����,�m5���6Odk< �knʳ��7w5גsV���f��T��'�,�aV��ꅰД�J���ZQ�a��_�0_��������<]8�C��k��m����3n�"{��2�Y�*˟2 �v,c��[M����{i��?IS%)�bzlm9�k{�S~�O�Y����{ooT���l�
~}$���e��L�PX?q�@��.5DAj��r��_��c��2&L��mI�Ɋ�^�SZ�E�X}B_�E�n����<Ͼ�0�p�I9|Гzn�>G��=A�宕_h�Fn{���"����8�Ba����w��f^��>$9�W�A&{�T���byMv-�Pv��%_�Z��9��9Ͻu�:�Z��Mv�2�TyТ�:2�Z\`�p!` ;kX1�Ȑ܈�;!�ȋoF��/{�~=9�i�ڴJ�{��#��ω���ܺ�D�K���#�V>�	 ���.��ʄa��N͆��T��lƶ�\+����?����Tz^^x����އW��"��"���1	��&OygWd��j�L��W�3^�r�dzV3��;������! h:N����g`ڑ5Rǽe�ޏ�W�����{)fNrRR\��-Ӓɕ����i'�U��XG!����DӬxm�;�VL[�n��y�4  ZD)5(�~,;-�ő��'�Y��/d��%6��v�l#T/�{���l#OPXXE'�PQ 5K����gI͆\[���b��`�J9�1��ͮ幌��Z����Y����A�|���lǁ�A�Pf��Hb+;��0��vNռ"��R�-H�HR���M|�;��dڤwZ83�a�cv��0�������`�*��w���T�Fajz�".I�${{+��M�x�c��Kvw�c�Ŵrg.�@}��9f�)��I��$�?�~�3=��Tn>.�ZFV0oM��U�����ջ�}�	���PfM�i�uf�0Xy��T�A���8XqC���>Ռh�������$!�%��V��(q��.V���yjv��E���ݶ��ƙ����7���4�=p��8���$�������ʗ�s����t�G���G�.M��O"{�1�'�J��X&�>�F�@��=]ˍ�<+}�#L��-��=�����FF�5��g���~D�ϤT�%��
x2�3�Ȯ�c��6����f@-��#��4��f����l��4!��Q��`�����L���X���-#@e��B�	鞘{{��x<�ۙ-5qD�F���dG߭������t�j������URקz�]�'�ǋ8d�s�7N&�t�8/3��@&S!��d	u����NF`ުs�΅�����@IDc#+3����hC*��CG�b����H?by��/���T�Y�x��1PN  �����|A��s{��Ʉ1��C�7�;/��s�Q���l'DR&f�nU�~�����.��}
��4�JV��\�vu���#�wz�D�������R7��r�I�v�h��_�Z�GAtL�^�y�|9��#�2��Ҹ�>�?�[��2V�^@j[�[�dh����J�@���Ci��F�)�,E<�)5/2IT?aUQ��L�g��u��kR�g�M���)�i*��P�' @lZ|����DT͝f�����T1v�+o������*��ޡ0�*�D
I7���юe��3E��kwvϏ�t��I��Q/Oh���d8�R~�� 7��u�v3Z�W��R2#>��`~��	^��a�g�Z/���$�l_���y�eۥ�d���dwZ(��C��~��y�9݉x&:*6�g�Cl�K�����j�l���P�(3v�\��W��t؏]�����f���l���V�%��?�0���(��%8���T���ҹJ�԰��{�b���=�Ȳ)^mMD�R���f�Έ����u�V�i/���� �W����^{;���a/$�t�N�E��qFm�ɿ�\~H����b��a����wp�;!�L��/�E���D5+��2Q��|D'������g(��d��u8�s��CKB�Yk�0���>�h�uY		n�2�g�Nɤ�D@=��ܸ��
�(C�M�:�sx���Z���+{�.����A�Q9{k�[؈�%$lw	�c�>Zxl[g��e���"����i�$1N�U���kYN�>]R���=¹�|;3�$g�6ϫ�e�a4&>���[��š���`�W�K�Ew�j}z��F_S����V����`\�Ix$R�i�cMgJ��Ek��
�a��k�U���lQM~�榁�J�Vy�5����JҴ�4��vd�mĚ�r���_�Z�1��q���:~=�DybA�f�`Jmi�*�v��p`��Ȇ&) ��V%��O����pqV)�,�k!!!=ʐ��/��ҞTr��s:sY��>���yN# �'�$sry3��^��@bi�W���5�`��4T�x��99;��Ϻ*�b��8���yzK&0֡S޸�6��d���/Aϣ�F:zj����M��)\ָ��2
h�}��n�ئ��|�!��_!�>_f[���ӊq�VՄ����D��������%�X0����ڿI}M(��ဳ��g��	�J�������E}�Z�M��=i�WM[!�|' ��]k�IC�\2���fわ*�I���mY+�)vg�_�`�99e)��e���!�d1?I�5c~~.�@��ɳ���	Q&p�n���{?T-�ŀǳ�����L25�I�8�Vr��W��ݑ��</3��Nu�n�I�c{�LH�荺L:���z1�`v��P����+��X5���Ǌ�	 ?\恳�S6��ů����@2�>�x�F���ӌ�j�4�<�''�,&놐r�X�7��׃��l�u[�Q>p���hu������Z� w�>�h��$=�K��+�g����|J�?��5�D�3��Hӛ~�κ�W��ڣ�Jg�������G>9��;a+O�OT2LH�{���&Ji
�ͲZ"C�i�ڋ�P�T��Z��e8���YM���'>Y�T�rZ+y*����'kG�9�bhh��p��ǺՊ!U�!VA
��X���RJ��m!P�fS�+�F	.�xQbs?����R�d�;,�@�`#�3�A�G�aQ"I�>M�&_g;����̕nc�덎�}z���un�R�M���/i����P�V�-��k9��V̵ц'�|�v�����=�|��8Qæt��� ���ޓ._.3�`K�_��v�Z�����>��;I��m��U62Y/e��<l�y>2���郜�vn\�.��SB�� @t�{��WE�8H�����U���P8$���h��`2��3�3�_���v�h��uw�����*�&vڴ%,�*9
���������*er�eY}��Ԁ�+uXjq�Y<��'f�=S��;�"tń�Q���n��;���JL�T�o�6�GR>Ӳv�?��
}�j{���;��O����ؘ�l�-l�h�z&��ϰ7n���nqŸ�:��?ܛ�v9�J	�S\�@"'��i��-q�b�^[I��<����N��v���ЦmG�l���j���+V�t�]Z�۟�@��}�C�=xuPC�r���?��oQR�&0��I��Az:-�35�=^z�գ�����k�33��g5�<*��9�l=�d�w��D��v�ָ�3k8�e�Do#��j<����:?Z���LMhE�#$8!��L(2�Ӆ���Ei�J;�W}��o��<^|�"5;'E�R3g�ªki�F��x�3 QE���o�M��O��c	O,�[��@5��V]��1`�M�����G���˘��>�Zb2j��xn��V�
}���2�&tZl�^��W�~��-�����N�ht9�'w��+�[�=��lTk@�����WE_PNo7u��x�y�Tz�r�,(�ћOr�����eJ���o%�䔲w�u�&\�'��:�S�P��6�f��k,�no�K�ݸ]��^q�D����p���n�������~A9+pt�🮩��������=N����3��4��X�3�9����/�W"+�H�Ke�o��i ��!�P��*4��a��K#�M������s�a�6[5��隺��qs1���3-�^��/r�(�4	�ќD������$P����nHF��NLM�b���֧[�E�[�V6�Qo�l�4���5�y>)ϡEbgtJ=DG��9���y��A�~縨�k�INw��D����3��"oPB�Lˁ�v9���5' ̯��N��~Y��Z �R��rT�`(�ڤK{�^�y�@�F�"L�$��Y�`����}������1t"�9��~����|Q����������7(�p!��v��P-0-R�/�wʶ��uL�/��q>�t�jY��G��_�����jO��(w8��'����OP��'1�)GwR�[�� o��Me\�'Yr�E���S
��tl�3��:�\�E����;O���������s1^��@�;�(����?�1��sDm�Ui%[�P��v  @�`�4� �1$Fo���cD����z��/��hͶ�J�Щ�d
�Y�����co��vX��u*�(�w��=yB�E}K���[4t��6#P�` ��,pޠjJOX�.�Y�Uqya�Tk���a�����<��m4�"�I�ʊ�l�����3��:�d����RJ�p������T/�F�?x���c�������q��/�Ύ�#�����bH�Q�O�<���3)�w����:X�w�Zn&-ys�ǞO�'�����$��Y��N3����zu	�c��̈́( �.+˧����A��2&g2����)�?��0�u�r��t����cW�&#��*�)�S�6�jUj~�'c|}R|��D���'�lS}�ڷ�/&l�-]W���,.�Z��['��ȪwJ�v���(i��25�d,#��=��`>�ݾ�ӶE�޷󖋝�=��?�~�8x�h&�2h�|R�$��E�[q}�e���=/hm̺�������M��Bc:�Dp��|��dgV#;�������	�%h�$���~f\������&�t�\M�S_�b=�p¬�l���kT�h�e�M�.�˛D4�O5I7�
`�g��!�۶C�	|���[�~*yF���5aϭJEr�zs�%e��bj�������å��E�:���}IN���ٙ����W��U<���vp
���Di���䘕���MN�R1��Bϭ,[_5̮�:W���q���z-�u�34瞅@@Վ;a|�*{���S0}Q����k���i67���&
�.ƞ#I���<!�c�~�=@R�ϭ���O¹�C�e��DX|�0)KHи~��ȢuQ���߽7U$��нF�3;;T�ݣ.?�])5����߲K8����m�ӟ����������gEs���sC���^�fwny+ɿ���V��H��eJ[֪Ӧ$���ϵ���_���;�W�vé�e���8H�T/i�/�|w�*?h�m�N�س4��n��;1��pg�tȧ��g�-����.k�5o�ɛ��d����2�/F������� ��|��	mTN�3���2�����o@��c]d����������M�'�&���r���g%U��\|xD�_DD��B���>��CD}o� <�t[a��2{2`W$��2W�v־�/�f&����w����Uc�����h5����0U�``��e?�ՒJ �	Z��.��Uf�������}�(���I�*Ŝ���h���mrxP�W����R��Rcj�|�A���c��On0�4��a<��!,���SܼHuc?�|h]�W^Ɩ�������+>���*��<�+�n�%��"˷G��&)�i��ΐT}m���@��E�J�I�C�ت�Y�����2�-��Z �l���������n|&�!夺`ł�@J�i������@�uwp��/�LOk��<�u,�4���ˑ��&+<��TdC�p�r ��5y�-���4���֟������#)ZH�C�a<=�]��}��̋����F�~�'6�ڛ�Hptш�C�	�� zqA:�|c�m��w��R��g�����S,\`�&�w�bmU��8�cb�U���)���6߆M�Y�'N�3��"U��tE����Ѕ���\�U��C�H����?3z��[�>i���	��C�iz�*�;a��IZ��a�*�`N�3�p
���<��z�$Șʨ��K,9N2wU�����ؠ���rS��L(d�<�EU9;�l��PRV�R�4ty9�L����%!uY��fUh�9�zQ}�=n ɚ�]��}�#P��5ެ�-m�O��7�>5]]`R�y�GE�����T���LQ��^ʃ�^���o��Q},D���{+��[���v9�6��6�5���]�5�_Zq����``�ח:��� FG�3�(i��e�+Aa���f�΅�}KbY+$$$H�̈+�<�����!��R�olL�T�\L�B���eԇ�w:�T6���
س���"m�A���x-�6��_���KrIZ�p��9�e=�E*�ȁ��{�%��z�T��c�r
v_GLl�� Ps6��*��O5�_H�ȹ�g��932��H|������_W
�iQĈ�om���:��;_^6��1��:�e�Ÿȏ#^Y`t�6m�jۥ�%)��L���u>����e�h�t�ƙ|���]�9��&n}���S�Iu�d\�W"���Z��v���������p�#ܴw�&(*�[�Ҁ��눍�����O���e|�Z��Dv&���!<���˴���;9'����3f>A��я4�z��x�$����9�N�a���*7�Sq�ϰN��~�/��C^$�R�ҝ{�3��tj!Kq�����T�n�n�j��r^��A�@롲+F����UR�.:�Wed?sr�mdb\��m�p�D'߬v�/{C�l+�Rv��X�X(/.$�5�7_�X�%�w���O)dxON:'���|02���7�kŭ�L�r��ӕ BO�4����h�{��A!߰xW䖛��`v.�?��Eע���q��p��C5ܽze��j[ �5�趿@5���@щu����{�9�58���,�8��_Y��C��ܸ�!x�rFH���P�r$H�u��� l3����x?V�c�wR���M�a���������i����}$���M9�!�����n
�6|*Q�����HXr,�_�_�dXQ�Hg ����p� �g2>tV�[qw����"�'�T/*˷�IW�}8��(�am،�6�
i�~½�1��U���^�}���m$�9��ӄ�x�r���Gz֑�jw��:��F��(PGg0���Ǖ�}��rۿX>Kh��t�O>��6�5H�q��]����i*�g��#�FA{{������g�o���/J����;�B����&��防|~�L�%L��Q������D�ݏ�y���;����ʒ����i�ՙR��«m��&S�n�K
{��=�棴�h�̟汗�F���-Y_�E�[����n���AΝk�҄i�q����c�y�v�ҷkP��u�o�+�md"�~��CUݬ
��[4Bw���m��W�Nl��Ś�J F4�E�*��4N�b���cW�ƍ�j�0K9Xe����Y�JNq�x;֭���fKǟ<��~��5s̒6y`6RO���D��m��ǂ����Zķ.cv�
+i�`&�[S�]~Ӝn1��1r!��t��kqQ�t$�e��������5�+����i���4*�I�q>�.+b��ئ-?��a��\v<��&��&�S��f�(rH!->��`�y�\ #-���z�{�eD�͐YUB8kl�v���<��{��
���Q
�4[�Zr:=�B�I��RX5���,0���J���)J��+�{&C�BW�$f��Ѻ�;�v�@0V��?�#秱R�9$��������s������ݙ<�Ǵfuu�H�hF��Ne��X�.N#I=��*�:T�k~}_U����G��Q\cSS��ҩ���$5� �����|�/���
1o�j��|�A������B�:��"!�N?����L��E+������,�QYO�AX������/���9�&PTg��v����z����}{(����4�j���(�\>��了��B�~ya.���F�=�L��x�I�g�-/U�k�FA A3�E�u/��<���ݨ���tOZ�]E���� ������L��JX��CQERI��$J�>woBnr�2!2��$�~��}�3��9r�tN�v$�����=�:yc.�̺G��iCp[1#2
���q&���<❿V����%zE��0�M�˽^X�w�#R3�)���O�.BI�&�'/���E�x4�B���5��呢H�H[v�	���9*�sJ'2�Q���{N;A뗚-�;�3s��,0O��q���� B��5�2bb��N��:�q�cQ�G2�sr<�Bߘ
l憶�tt������=�\��������/���%IZ<Kl9�q��	w	 �������4̫��.���n�/��L��<lOq�b��^���[s��F����n��<�U�0d�;��0<�i3K-�I�.��f������E �5�y����M�-�GFb�@I��ՙ��$��B��F�h��|�4�d{�kg��#hj�I��Fzhb~��d���a�)�Z��X����&>b\��U���s˷��Y��ae$���_�����~�o���/�O�64p���Ao^���-h/���D�E��$W3�q����qA�۬q<�y�(͘�)#��������v6I�}������o�=�~� J�O���T6�1 �~��gO���t����Ƣ-�XH��i%+V�U�'(��׫��=��-4^.��i4S�l�o��}��Q��D�"]�e���J ����֧li_��m8a[�C0<*��3Ы�z��]i���Y���'
�9��S1a{�dqvчea���(0����ˉ9"Kʽ�5�b����3����׬�ɛs��Qj��DqHD��^[�
Sۧ��Y��衝s0ǃ��Q����B���h��/�?;��ɤ:T�
f;z�n����2�\��
<P	��i%p�t��#Q]� ��9P1_�RG��g�z��Wve���*w���3���b�[ey$\�l6[�s�x�M���Մ H���=�������/﹉������``�\]]%����!��!���1C��8�Y��|����5G��Fa�V-��)��p_{q�US(��y�j;8o�&�܂�2߆!u ����{���tg2�bH��/q��L�sȭ�.��";�4j�N�516,�����}�⼄t�My֜��ۣe�Ԙ�c���I�e�2t{��S�/#7�'��G���zKa���dz�z jB?ԿpZ�<|���
����dq��b�3��3K�WgJ�!l����95h�j\�I擄�˰v�� �a��o�,��x妲x])��m�og��)�{��(�� X�T<	V���{b?��xB/!~���N&3�ƾ����w}������mv�س��,*�&�YY6��`c_[�΄��t�m|�ĕ�Q���#��.yPx~?E�hZ��`�{+¬nn�e������]H������]����Bd�ko��8U ��0�5;�F�77��k��e=����g�� ���=e��-�g�juB緽ПGD�+Nh�S9W�g��V�i�w�[35�%Y��g@
!/����[�Ȉ�R�ս����m�ـR/��X���9��`��n'�!�_�|�	�pF�tq��`('��M�B�|��A������q��ym���6?���˸�`Ib��6��i��[)��~ڇ�~A�&���7+p��.G_��;�aY�q< �{�<��ܖ{pR\��EÆ&
IɎL��.���M���gjڡǉ~L���#��'�פ$>]	5�*DF	Û� ��Ҏ�Ӎ!��� dn"Ƅ3�]� �Dѷ߱hr��G�Kd	]ޑ����R�Hܰ�3���q�_��6As(��)��p��܁DA@�5IC�ɺ���ƽ��
�xr���
TXĎ�i���a��1x��e@n,M�p�A���} ���I��EF$�3�b�@�=(�u���Ҏ���'"�WU`�}?�#L׉Y.wr��Yl�����i���
o�<�I`��xQ�vl�:�G�����?'h���f)ή���}�1�	���ٞI����E��4kLw^�ʕ����n�Csɤ
�0=�$C�\�oŪ�u��]�����'��~�t͈�1:�'�]�^Z�XV�=�c{�����|r�=�[�󄮊��u��X�>b�~�:�b���s�I��'q�m&�)�W�s����{�1|a&�V��H��ی�n.�3�����A��^�k=��C�tePm�0���5���u��Y�LsHc���� a�V�z%�~i�����Y����BT�J��2��s(����̽�&�=�[&7�=�n"�~J�W=�HىI.W����(a�Z�[�?O ����4\eX���FA�AB$���;��;���������Q��ex������}�<gN�sf��,����IL��OR�߿��(�I�����**V.d��x������0�=[�+#�0�jd��m��f�W/~�ځ��u^g��:��L��H�ј>�tf��n;8X8���%cO"hꘉ�x-9?�<h�R��hN:?ۻ�4�$�I�\ ��f�։���\ ��~]ڑ_cO�{w�8��䴭4%G�`���'
���忨�@����Q���(2i�!ʁװ��u���6b�@�e,#%����x%Α% z.��6i���V·�gͿ�L�Y���B���Π�跂����^�g<�ߩ;�X&R�3na�l�=��O7.mj�[�������t�*_I�m^�bXW��>����Ҹ'���mS�v��C���<.�mh$I-�%�?տ4�"X*N4�1Z��5�h͗-l7�G)��
���ޖݎ��L�&_�lQz��CB ��F�R=�<��3&�4����t�خ�,Cn4����#�Y�h8X���B�Şm�i]������0_���V�I��q6�)
I�Vy�A	�[Yo�U�l�T��;�����p�e�)l6ԐB����eЧ�"�^j����h�P��h隿Rd<N�3#y����o ���E��u������.�E�-����O�5  ����)�S��͟����?��\������[/|��� :��?1�"�l�ܓ��]��I�E|"# l7ݝ9��	������ۊw̃�f��;�.��@E�`�����'�\���:g�L ��Q���0�Q��P//}\ט�_���1�a���!��^����P2�m�j��U?�OsM���ݳ��d�ji?�N����&�E�7T�֠���e=2jo�r OB�"k��#X����Ul����%�ey�	���#��``�j����dH��R��4<]x�fʰY�)�ٹ�Bf�M���O?�5�!��X2���i�''~��	)�NH/�����#��Cp}�H�Y��PkE��U��$�`9��W���܄u��yO\U�������Θl����CN�l{�N��vk}�jQ��')<�hj��_[L�*�;Zx����;����r
�����\���Z�"��%	7oH�u���g�F�E�"k{=�I!���/���+ [
	G'�L���l�Z��}�!��>�Z�&[����#�������H�dQ/-P�# e\���5]�e7����@��pܜ y������u��aឧ�&��82|�ʉj�1j(G�S�yp,7黣q
�vBmh[���Rb���C9/������w��0�<lt���+A�LIy�k���Xg���<X��ߒŞ(b-d'q�M�HV�uw׌��f$���D�hld̶`ws�A�@���vH�o<�K����1��־����R��)l�+����A
R������ν���K��I������Re�{���5���،:��#M*C._�ψ���f$�
g֨�	�������L�=�V,7�\��уJ΀�_v:C�S��ڐf�Y�}�[G���｣g�3tZq+�{dX1�=(�(A�zRiI}�P�`�!k5{�k)�ҐՒn�CI��s*3�÷9Y ��o�/oTX�����ĭ�u�w�~۾��+4@ ����{�4�
����Z��h�[�M�"fUZ���;�z��-|Eŀ./�L:�uˬ�sX>�`���!
���7Jb��2�g�3,
V&��B��v�B��0�QF�y�]CB��bvی4�@�N7`	��fdJ���f�yc�U��cHx�IYo�r6S�G1E� �EΛ�߰Y-1���f��X������ô�����ě0d�9J}���vl�v
?���S�nok~P�;�ɚ|O
��)0����E8�wh������W��_���vt�_������W�?����J>�!��m��CD���}�{q��֮��i�l�hÁ`�&~J���!Sh��I�F����A��nq�9�3��;�q2m����̻�A*�Ն=�!�����9_�-���Zub�t��'��-��*����̃��;�X�n7�X�J�峑���#��J�N��t�'��߬�0��oP8�ަ��boh�ޒ)�G?��+J�Ls~��9��[Ŧ�,$��5k<��\~������j������ϙ���K��%Cb��xyu2}�� ����Yod```v��[���#H�V��u��H��t<�������ho�R;��� ��_������]@�+�>�$Z��Fr���·0��F�<G~�V��G6�QQ0"w�5;��d�U�/�R�,�r<aܾC����)!1�D����k$���E��7hQ�o65����n����P�V�_"�C˂�>>֋�[�{�(g?�6�a~��1��1�WG���7|�?OF@-,F��$���a�PO�!U����~_Fxa�%��Z��ϭ�ԯcZ����"kDB��F,E���������k�wb0��Lb)'�8��_��
��&��w��P�Y�*��l)H%����������ֱ�0~bd`��a�{��OYv�����f�_��@��Hi��Ú(��Go��ёq�i⠪$�I"��Hu]�H}�t^�;Z[[���*#�mM|�"�:+Ӧˢ��&栬�8�xX����JW)�o��@�/�Ѭ���M���^Y�u-��Қ�UPk�2Is�[�2gZM�47:H��c�JR��!W���a���� I��^_��թ`W/א�^��,����K���Z��]�K�#H�W�����j]��Q֦�~p�Pt�[��W��A����3p� قZ�^���QR�(g����r����������a¤F����<Tm��_���m�z25�f̓oMʏ�D|�4��pXcy��1`�L�.&�:�X�����k_�:�ٻ�-\�lvoe�p_6\� в�¾I�bO���g��1�rɛ󑨾���Ce?�E��7�ą�g���Q���\4ڣ� �+�׍= �ZRX=/��,~b��>�EnN\0����e|_����8��jQO�XVzO��q�%Y b��T�F�d�����ax�4���L�#�&c�^��U��^A�e`���2Ν\ٰ�$|uh��l�)q i4I3?_4Sn�,���(#��׃C��p�o
!�5$(�n����Tٚ%��.n���'��0`i�0N^�/���-:9Y�m����l�(��Ak�^���dKק�-��[)sP�V]3�2�l��"~�Gb9Ӎ�H�
8H�/�ū"+�#ʯ�R�8u�n�φ�JK��i�1����T4#,	*�+|�������}9w���NwH��}JmX��C$�~�S���b]Wꥧlfl��󰻐��������QT�	2���?O�K��#�?��!�{W �#�����5�f�z���T_�� ;L����>$:�C�w�T(k]�ޗ�x ��M���&�Op�f����/���� %.M5�ʬ_P�ăF�6��<S+��`�Q�9��������e}���Y:����%��J�GB��xN6���T�|	z��ԙ��_K����I�n�F��r�}n�*@�X����B&���9髬�P̑*�u�f^��n���-��@0/�#̉��9L�s�Y�v���mho���Z��T��B|�*��oR�_��0m>A����H��@??���������1\�2�N^�@]y �Bjm�<]=���l�h���u���V�W�Bhw�h��:���*��QD��&�xj����c�e|��\/�K�O�œ�BTp��~��\#���-���L�̫Y�M�-�s�7�;L�,+��mFT�p]��{�5͟%��Ђ	)��`f/��"o�kp�������p��(�<���3�r��;7��;��
vu@�	=�;���-�P�[@�����7�	0p��׷�1?A�a����Ĉ'��������jEP���%_�D$��ø�Z#D�n�
ǌ�Qө-P]������K:��������	a�����iP�3��%_��w�[2��zG��,��4�W����Z�g�uZ���u�B-����8���BЏF����V�C�Z6��#��;s$�� -��j�ϺHͦ�����jQ�!���8?���5�w�#��-���!�;�❄�f �ij��VA��{��ͽS�EVm�2NQ�JeZ���Q$e
u�$.�v�=�;�=�W��?�F��{�<�)#�̔e3&�E+
�[�{��W���yj3��9Q��7ˠD5XQ�8�3Wd�Q�@E���I�<,�})o�s��U��Q��װZ{�gUJ��E�j�W=��p�s��Z{�[�:\f��裄N�ܤ�� ſ��m?|���_3��,U��kF$�*�� GdJ�##^�v{��[8�[ig2/���D���t���l�P�e�6�S܉8g�+�DO:�7a��̸|G*$�~C&F<��a�ω&d��v�V��V�L�k9`�C��d"�q&s��_��|�~�iv�e|��`MA�#;s�T���V��!.,��p��J(�V����J�"-j�+0�-(�L&�T��A �O�ԴT��&Tg�F!����EV����f���Sh��F�����"��!�᳼ro��\���F[����D���̑c3�+H��*?T����� ��%¸�d
&^Q���j�j��y���%�8t�݃n�5h�IR̷�צJU��^/AǇa�/�a���ҐX,�����5��h��j
ѿ��t���fRh@�V������`���[����:x�#�/B�yߥ��]�1+��ǲb�gO�׿��'�z�ێ�D���Gh@����tݦב<*����`�h��,'q�W��Oz���	�d�U�R�"�}@ߵ����w��{=����Z߾�b�P����9���Zf&�����+��C���ˁ�͓�=Q� ���W�h��fU�U���H�s�	�o[[�I!9�v3 �,dŵ�%]�|{�����y�a�+�c�Y�֦�0���|����B���|,ƭ�>�A$>=�=����E2�, �1)q֝T�Yn����`ѲL|��'wW`E'���� ��!06�l��˲�z�U�?9Xٳ�sF�q��5w�7T�D�V�D��/˿� ,C>������<��аQ�&4�K�U:�$^&?���nm��8������~kɭk�1C,QDT;�����]�)tk�R�*Ne��kF����/J�p.��)�O���m�L���"�����eLxS����^.S@�t��A}�D�&`�:�ն��$�b��íQ�yHY����5:8A�!�Sg��qm��/��S��t�U3����Zx��m���v���@4��n��Sl�ܹ��	*�C�!�ԁ�����:B�E*'늆�W��q� W,u�����j�����W�T��v���4�9/
�LEj�0#���S��7#+�ޒ��|"��ȸBD/���fAK�.Xmߣ̤O83��]o�jk����#���d&�E�k������[I\�T2�>k8��)ڦq�4��X5e"h��v16�LP��[=6�Ds�=Lm�PwҖ �X���-��Uft���/��b">~����X�,�	�L�~g� ʧ�	=։O0���'�����f�b���������Y���U(f���Sj�JQM7��"�0��B�����u���?&�g��3����c�{��o� *�n�0\��3�w\;��v�e+Jyfd�To�C�8��D_1�_4i���0��q�İ�Rm���);��=&���1FX��(��f�g���h���|]�@�&��$6VX��
���M��g�j����6r���P�ϥ�?��q(�� ]QE%n{�6�A�I���jU��s�@k��tC���h��RF;%S�!'��g�Wl�Pi�'^��͠K�āS�"���Gq�u�����T$o��6�2���&U�!hW��e��M��R�r�P���lpFk�{N{>Y�*�L-�U����P���˽>9�$�6W=ш�&;�W"���K�f)�* ��³���Ջ�y�	��Q��k�����'\�{~��.�dXY-�R	����%��Boۯ/����vI�CA���r�0�%g� ���bA�i��K2n�qƼ,ƻj=��[i��G�'�4 %e�b��4?E"��&�����e�.�ƚ�h�`�XU��@]���w}���"��m�G'�s�t���S�׌�yn�P��p�6�������D!9Us���3{�J�d�R;1�]���gN�*#u;K��(~S��`�Cf`ý��V$짶E�T�u���IHd���;��fn�gV���Hd��/��O�v����_�lڇz�(���
r�L�
�o���֖˪c8�7�}�(����C���m+�DƦ�)`k>�ۜ)Un�霕j��1��8��W/_z�H�N��jU��v�<�Bw{�Vv*1j�[��dvĈd����09���ﺩ:`�Nv9�$AK=n�/R�L�5��,h�c{��8�����<MT�0��\�س�w���6������O�s.��������F�,�l�����3�3R6!��i��D��g3l|�N|���f��#�i?�c�x��
V����Wsf��X����"+��a7���;���5M�f)��C=)�$r|c��靝>�������|b]�����\a�f���vj]�z��6JrH.�jk��z�χq?<l���S��NA�/�Qj�!�����?�0̵��#hzc�s����HU�Xfahui�_[���7N��ͽ�fR������ZM�)*ҭ���q�H OԜy6��\?��O[�C��B��Q��i]�p�fd%�1���G��C���4�&ƀ���u=����5��ڷ���*f�ꏜ��[��֗���;����v�R6�ml�?�e�f�׼�h����0�6�h�~�>G5#V��ʀ�&���%4�Gz�o5yzԻ�z#��OaE�H(ע,���a~�kOq,�]0�*3~(����9��v�
����\�|�k�8�<cp��l	����n��C4RO�|��]
)1��UY����3iH�1}IIZQ��NU���Nn)�p��2��"(�ӫ!(�
>$�=��V9���Xd)v���X����<&��U�Q����DH��/qjo�|��S��/�`{T����	��ʈ9�H`�9 Y�i�+x�l��+Xv;䃆��-��D<9�ϚthY�7j���H�]��:-oh������Hh��4=8���j����b����t̂f�ĥ+��~Aq5_�N;��@���]Z�-7Cl�������U�@n�o���j6��+�ɂ������&��g^��<�J~���D��#����OѾ�-w�Ql��_������!f�纭�ŀ��9���^�Ʋ땁.�~��K.�/�`��kި[�'ۓ�v�c��������������NL��7�m����߱��ZfFsg:t6>>o� � Fa�ŚK���=�v�#��d×�xf�]��:��p�N�p(zpw��o֡@ꔺ*h��T$J��kOp����]8�CQG}��i���|$E|?��77%����=|�����Z?m���\X�z�y������~�!�,�"���S{(
	��vQ�׵�^m���Z��ƗC�o��R_�-��N��㳪�9��q}F��6���=G�6�N��o��A���g�ݘ��;z8��+��#?����ZH��*��6�)%��8�y×���%A��FH�`S,a�,�8L��>Ƶ���"d��8���\������g=$����w�"g]qhȩ���=�L�T�t�9v�V����8�]�֫^�����/�E��W�KDFH�W4���M>�� ?�ʁV]x����,R䒞9�	��T,�̿ '��z��=߅���VES-8�z�v�:�9CQ�}T�UC߷@��Y|�5�R\��6Z��=E�&�ʪ��.%�{�1%c%��JS/����)�Ǥ?.c��՜؉W�3�PnjQ���Y��z�>s
*��XU!�X:@�H��aikT
��%��U������%��F���EA���׀\áhx�3P񺿞��D�#ғo2�U� ܪ"��O��
�w~�����e穑��F̑��̸��l�&$�΁]w��X�a�cR�m;�:�K��pv��{.�y���F�GY��c���Au��d-�C+Vt�U���W'c�L�t�ܠ�O��l���jp�e�B�F���L�1�ǽ�����qp-݆02��� 9�Qq�2����5��Pp�nyb�!�nOg�B?��IdU�b!�5_F�f�`KWS޶)�}T���nl�L�H�z��P�yB������$=~��J�¼Y�m�򷌲�4���pτ^�6�|f��$Y4p�P�Cq�'Z>wĥ3_��sZ��	��5��G��H��Zy�$�@oJ)�ɓ��7*Ǧζ�Đ}y�Z�%��8g��ь�ĕ���?��y��������e�>�$��|q�E����5+8�8Lbb�4�H<|eAG*b����_�6K���ک��rQ����j��~LJ�s���#*�S���
���EW�E	Ne�ڿS ����Y�gm���WED[��@6�e7�k��5��氬��YQ���1����n�a*P۟D��P�9+v���4�W�n�cƳ/ylpE�Aƛ��P��O}g�7&��z������W:�M>C�$�p\ݝz+X�S�v��4����0'9���&��M�i��G�)8M4r����9y�K��$�tSO-���|t\�Fa:����<���a|Yl4�i'���!l�lh)<Ȧ�G�?I*��E�����j�uvqQ�ԃpO�7v��~cn�Aݪ�ǵ@%��@&���Ӝ�\��)#g�P��x���o�ą �ek��t}�Z?��Jc��tь���c�c�s��Ȍ��#���3�Z_��n[M~���a�~�")M�K	���s���g8����y`����&e�aEB���Z�α�
ݜ��c��6Lp������g��Ns�ʳ���䗰���N+��W�Cχ�m�蕈�C	]So�3���l��a�ǣ�f��<�zCm�"I���Js����~&ݶ�=վ%��5��T�/f m�S�Bl��El
JS_���d~c�9ts�����̳�Eo�j��L���ƭ�H��[<��fDU�-����pn�`�ZW��TO�Փ����_�nXre��)D�v7+֒�ʅP_��D�O�'��]�����6#8EK+���S��qt�$�FwKr4"��2���x�vEK�>��tww_�z����w��a�e�T�g���9�yVI�h_a���;�ш#s�"�7�Kܞa��PRD1����TOLԮ�a��N���C�r���^I���]�dJ��Bd�ݬ�r�Yi@?�h���$F�yg�ק3,�aMP��k�m��|�3J�F��k3�ń:�{(�/"<.��A�����5�:�<��������merZ�����\�m4W1G'�m��Y ����s�b��2
e�1�a�NM�s���d��i.�Gʴ W������V~j��R�N�f�5�����E7����_Vk��O�65�̐��]�NXҚ��aP�4Va�F褰9�%7]zڝƎGdɐ�*]z��}g³D�ڟڼ��xѼ��4� �oҡ)h�~"2@U���t��m��G�I�����tbK��k
�!$H�V��62�h�t�dm_O_\Qr�� ���Ɖ�U�r����Z>4B3��n���n�}=�6��$W�n���ԇ�1RI֒/l�c�8ş�~�8���Ґ��:�BzIv �榆��c�Ⱥ��{O���C.�O�L��JqZ@�
�RV#��}���b/�J��Uh���NL��L�M�{�u�q���F�\I�01U�*��b��9����!��&�W�X�#�4�P޴g~�@��ژ����Yf�O�X�}�b��_Uԭ,���@W���N�����;�Hf��a�P��piZ��2���nD#���An�n�a�į��X86���fB��]J`�.��bt�2[s9诿�����Зpyļ[���BA�8�jқF!w|�3H�J���۪'���Ń�l��
L�,���z�R
�D�B�W�6	O��<f�R��^Q���M�{w��&@F�&G�C����x#S&n�ꏍuɎ�PÝ�4�uS�HW���[����S�a�z�d����E>b3e�v5�"�fK��ߥ��4�������5n�|A��=�Q0ǦE�pߛ�^��,�ԕ����*��6�#:ήQҴ{ǰB�k;���&�����8�܈��B�ϕ35I�FH��a��#�woZ�?4���������;�o����P3BG�U�ϐ�TI��1,���2Ӭ&S��F/����۸�u2�������S��0�,P��.}u�|b@+<|bp+���}�ފ8� `2���A
Z:�5��H5��6�!ܵ��(��!���;*K�&S�r���������c��䞩�
�7e�XN�Y6u�cxi�H�Q@~�ɫ̌��Yٶ���A�P����$� ՜R���X�Y���nM�b�͌��rt�)��bϔ��bӓͶR�[��C���[.��lƊ�l�?9(���A"���JD�-%�Rw1щ��YU��U� �|2y�u/���=�g�%��4p�g�$;ƛ��q�6�϶5ٽX�T^�;ҹ��#���`~�*,a���e8o!|d��k�q6�In�Td@���?��5F�6���vN��ͅ鿙�Id"Jh5��c���W��*�dɶ��SР�����*�5Z	�m�Җu�3*c+Z��,��ˠBHʹ��s%�͏�k��ꔜՒo�t�~�R��cn놫�.���:.഼�a~��kG ����+�������?t��!��$��Lg��*w����#c�:E�j/��*��[�ͻ�Pe5����&��?�J�if�T*�����{���7(B��GT�a�8�A����p p�q��u���sڅ���h(��މ���f|S���s)��{`^Q���D�:�Q3�m9�_�c�X��K�ڔ��� �
�U2v�$}�b�	d�#6E�o �3rP�"��6M-Y���n$��7H-�S��/ӣ��|o��=�o����ّq
"��V�5�i��)���e��f��XjTg ��+Z�[�IJ}��J6��P��@��&����X�4I��D�O#q,{�9��s6�̽����c92i5�y�_����@�6�H���B�5�[F���_�t<��C5�N����3�l�N��Hc��9�(8m�*7�Cv����ic�j��:���𬚻�Q����H>��k�y�}xm�
�S��Om�͛�܋1����Y3���,3�I_�3���>�IyO��BD�����맖�1Gзj�������,IZf2	N5�p�ߦ��p�9�X5r��d�U�-���?N/	r/���@��o���&f����k���L||����ᢧG<F�w�m^���.E攺ߺ}��o܂.��:���,�Ssg�#��@u�	����0=Z���:�گk](IU��k��H���b��,��٠i	*<��t¶���U:��!y��l�m�E��RD��:d�^����8��$��{��0�P�͍�O__]h����W<��;;��p�e9ت��]�^�+����޾���R�>��Ra�;�~�Q����/�2��|��f[��瓠�:�o��a+433}Z/7M/�OcCJ�KШm���k0#�Q�7,	�-��MY	g&B]�m�� �P>�����I�Դ{󇄗�:�'�p�F�E����{��ojžr���.���Gpp�ǹL[��q�2�XjK�H�_�Xm]_�Ŀh?��A�^�NW���O>��>�ĉ��V��%�|�dc,y��K�!AzU��Է�/+3���Y���۫px��x9�fL-_/Y�{�xh{�ۮt콗�lz@I8�#^z����k4H���L=q������Ͻ;0e�?X+��q�Б��r%�,����r�].Vx(�fM2���{�>x�z �H�[������ϼlA�O�7&�͊�;ދ�Qw����tu|�*�tV=Xͽs�
?aȪ���}�]�p,UZ�bj˵Vj�ת15ޝ��%�A�k��^�3�-GE��i�E�i��sQ��Ӷ�K�C��M������l|4X��e�������a��t�A�ś͌�Qɫ �/����s���_OH_v6ڧ��_d�� ��/w��!x��cl�RЁ�?z��V/՘���2#�u/���$��݀7/���9�!X�lKSS�'��'���M���|#ŵ�I����Eb��%�\��mW�3��<P��婧>�=r����:�����)�P$��pu{�Vz9������z7�_���ޑE��	��L���������_=��'/�~$eROi�3�E��ej�u^V^�{Ɠ"r�H����^��n�o��N��c�;G%ID��R��N�O�*�ӟ��g��}���������Ӷ�e���-ƒc�K^��3�s��P��
]n����j�෕z��tخ��F�
��竗&��`җ���=��p��@ʂ�-Q�7��Ғ�ǅ�P�NW���k�cr�c8DN��9
����M�׍��ٺ{������뻩i�ǻ���麘Mc��A[���U���T�\�B[��#�� �N����d&gt*��N�*!��|����/�M7�L��U��b��	�"2�r7�ӧX���:K]ϝnˮJ7�c�J?K�fMa�E���}Y���d���̅�@�k����3�\U��K�E)��/i��6Y��ˣ��ֵRʦ�I���,�s<H m��꺺' =--鋾�^o����!/�Ew�U�S�}�6�?��`�*6��ۭ��	��b��ŮHKo!_��:�Ѕ�l͇��=��%T3�d���Q�V�Ī�B��f�(��9; 2����r�� �N¶I����rR'��R���9G�J��|x`�5|1������h�;f�=Y�ߎFVVs��u�$|]����բ�W.��Rb�e�kΖ�p�qK�=��҂��r_l=0��w�����E��"hT6������7'��&�pr�-W���߭�����M������v���Qv0���%�S�|� � ����0���FJ>g-iZ\�57���%ۧ�ǋ2��M����5�I�������8�����H����C~Z�n��!#d�#��*λ�d �s/I�hVC���Kq��b����2����
x�D ��v��>�6��w]Յ�.��V.���y}�QK�S�E[�s^E}u��w��{F/�<&��� �O�}x
Rd�t7y8
	����m+��-Be�gz|�s�s?I���<��-�T��?�(P�"ʹ�~vp������B ?��w��9�O\�kXF =�4�þ�g�ʸ�i������u?�6d#l�y��2���ݭ��X�v�6°�u�aU���+��vG=�KY�yf�&bD�G����p1!*t.3�E�¯^n^�q�Z���|��zS/���<C�sEv�:N�^��+��+33
F��QkT+y�e�s���da�m����߿�1J^�o�.�\�;���I)��e0�u�B�|.��Hn������X	�,P6����M����1*���y�|K8�F\ե&)���lOc��km��|��A�)C��-���y�%>�����%�#~?�*pP�fh������f8P�{������*J�x�쇠X?S̾���{��HS+�N�d���'�n��O v!l.���@я��J��'�r�4S=yd`{X��0Vb��9V(,�b�v0�$�Q�a�H��������ޠ�\���$���������Q�.r�H�`^|X+7So"�7�&�Q+�V�����������܆ϱ���� ��(�ֆ�䱝Ehz���V��׍��Z��[^e'�,���榆�_�z [>����䔼��\㸟O<�n��V��zu��<���,�$�w���P�c���0W6�s�(r+�.�Ӯelt8�X�8ɸ�Cs�coi�����ҧ�g`�zqf�{�q���|48�T��_6ehML{{Y��/
oQX.@�_?�l�LWQ���<����]���!`�����J��C�Z, �{P+����Q�i����p�L��+�&���[�`4n�a��x�џ���p�gS����,�&�*����T#a��č��s}�R,�������ٿ2��,-*�G^b$��஘	��$р���TM�_cw��e���f5߃����Vb���*=��iox+�f9�����\u�� �\/*�\���|ꟑ~ߌh_��ϰ�Qm	�+��KUy���iX���N=�d�6VG�He/-��L����3�n��e�`�V8S��AA�A�eݑcbp��Ҙ9���)��ElX.?���P^�@�6���$�w�;������������w�S� 2��\.2�+/�,�/����
��g��d�{�J�+�������v�K=P���~�1	�=�Yx�e�B8��S�z�°�h����k`���'n��4OF��O$��NPm���Ŏ�k�!?�RI�fߨ|.,����T���i���������I4s�J�D��|;[.��<c�F�g`��Q����:���q�	,A���X�Q�ߗ\^�/�~��I^MD�^+���m�j��}r�8O^[-s>B�0��������������)]��$�ڹ��&����`������}^t��4���+���'��ģ�����<�$�P���܉~�l0Cp���y�a�T��:/{�Lc�#�u%wf�#N <*hwT��߅϶H �{9;o�����X�����a͍���l��+��4�wm}�}��:��,�I}Og�=����=O�3��^�&0��l�i��k�qoyRX�;���t���ۼ%�t�e�u,����� ��[,i�H��V�z5��w��0��`�#N.f��c�L:�-���v�֏d[*��;���w�7(,Mnj���Lxk��e���p/�y��Ӌ����D[.��ء����4uy�Fl�{H������թÏd!6˱�M��a�`A��rֿ|���n�)��g������
H�<E]���O��e^7aG�Q��r�u��LYD�_*\�b������t��w�F���������@��I]�Y���+��pέҟ�2�jڶ
ϻf�ho;�����72��<_O0/=l�<{��%�f��d�:�YR<�8�p=��V\+���SF~VV���s�&��/Gt��~��L��1Hl[j�T#�����,��n4$m����D����VJ;9��]qvj��4��,k&��*��1@̠�,��=/�7����w�'�s�k�?���[�f����ol������/�gb�B7~\T�2���,Ҷ�b��:ʫ��	���y�ow�-/-����6r�#�G'aܕ�@՛%H�a�>-լ'}:�������q��������l���_��W]��f�'��V�V��+O�,s�A�ά�[3I�+s�$�?_���=�Yܩd��e�W�-�r�U�J�d�G�6�]��Ƥ��;pFU{�r��QW��X�F�
'�G(o4���_��1�d��3:ꋫɄ[��V$=ׄ)��>ͨ2:�giv!�SůS�L/�.��L�b���\zO�:�޿Y���fv�� �;�u��(�\4����~��������o�r���1���ݡ���=�����t����<���{G������ƌ�	��� ����⨼i�d�e[�6O���A/���&'���S.O��a�R!!�ܾ�0"e��m@�V�<����dSZ�ٲ}烗5D��2N_㕇��s�fg[hV�f�WI1�0Zi���H�9y�(���+�4R�:i��q}d8kv���N�˚���k�wi�������Û
v��U�+�xs�>��o���T���gm���
rqSw����<��rl��D�cY��DuzcŊ�#�:��}���JL*��q>8��	;���.9^(��n�>,�p@�D[H�72�Y�ؙ���Y�J]O*�*�/�>u��w��������!@Tj�v+tN�r���c|V���!�x�ɲ�J����K�9#���T^yX��Ȓ���٩�P���P��}]���9u��ꦏB��
��P���	�����`B{j�%��n-��+��-՜9�d�'.�C=*i���8w��OW���QQD`��.����n�n����a����n�Z^���ݏ��{b��33g΢pWo�ԵL	�I�ظ%}]��ݽ�✦'����a=�'�UW�垻X6_��Ie	Fu���}H��Έ�����'*s�-!�#��k%׍�Y��Os�W�KW������4cR��p���GS�^�	-6��(�1�")'2k�S5������4��X7��Tv\�<R,$�� ��[F�1��]t�v)ҟH���,߹��Z����xrWx�U�1���c|�� I"���_�����c͋��K9����gvyV��#0>��s��[6�ɛ����ag茤{��+�s�7��Crˬบ%��X�jB��-��Jz_�������2M��;�I�n�Hf��B4�<�I!E�}oT���r�@�~C,����Ť;�a��Ӕs�x��)�)�3%%m�A�.Sj���^��{���HM�6��v>�~e�S�P!�u����N��H�����������+���7+L�E�J��#���]�zFb�<m�>a�󨍗"s���D_Ps�8�F�e+ɗq��~�[���&	̿���Re��Qz9�I'���u�AI�����y����H�����Zƻ�����[5�@����.G��ى�������L^�}����E߇ϻw#������#$o���_/�t_ֱ'����|-�A�^o��HѪ'�BW�3��H<�ɛ�{S� ,�hS�D�n�&6�t_�;���+ͩV��*��~�6!F�m�z�҂�X�2)2�S�v߲�:�_YA:5�\[/�_̽Ȗ�D�!����5�v�g5|6�WĄ���da-F�F>_������p @�
�L�|��d?+���/�[)e@<\Ce�Κ���cZ�J�u�W���/���0-]�w��q�Na�9�����zw�AMrq8���d�Ē����y�.��'f����:�W�ě��h�e]/.d��%��¥a$}R�Z+��E�_�c�ሦ�˼^(r��m�_��>M����#0}hH�yzr�d1#�s���C�?ٱ��(�K&���%l��Yw��
�rOK���k�&������Z7��M���.{m��|�𬓫ugrx����v��Vy��"x�Ԙ��t+�sݔ�֐3M)����iɟS�)�1W��/�5L�ϯF�]�V0�BL>Е�3�%Gw��q��@�V���-�����4�κ�;�|y����3�olcQ��h�	z���C]��e�i��s;ZY �0m
+S]!�a҅D7��~���5�ـP-�)l�kt���ylP���;���x�w��hN�Il�4���1�������c#<V��z��t}pQM��>A�]���a��_G�ѭ�n1l`�"..�L���g����b���2Cǳ�tf�}V�b���iZ�MUŨ8u����f`\Qk��Ȅfe(f[�ڰְ5�E��f��~�t)[�c-������>LE�{$�(�M�'������8�,�O�=]j����S� �3x$��I�Cr��������c����@u�N�x��@�h�K�~�.d�����O<�w$���?��3t���Y���Mx�`�S�ꏉ�\��\>/�NG�߳�=��*A4$wL<K'';��$U���G*�fGv�.҇�d.;��/��K�,�n��ehQ��F����3���<���<�A���"o��H/�4#.3�	��FDk/�}���]�#�3�ڪ� ]~��+)4"�%F��唭{,�eG�h��x�ql%�@
Ż����e��q�>��A�y/�Cǘׄ�(V�����#M&ǙWBտ�P�2`�e��5$��l��_�0]v�ڴ��]��ܘ�`F[�C�/Ϭ�s�{,kj��K˨�T���?�_��~��.�y���7���E_�r���_�bp��`8]��4���&w��n�u&�CŨW�h�"��Ԕ##U�_�1�Z�U��6�X>�z7�T{�"t���ev/�9������? ��k`iB )8�TtiH�9��5�?����N3V]���9$#��L"&���~��',���gK�A�o9r�l-T��Yj���&�>��$�Ft<z��
��Y�/j���ѕ#yY`!���+UC球��9q5��\}��i��R��w4A�cܟl$�v ^R�D�B�_1��O�ྯ3�bU��Ŏ���ꁾhR��M����� ���Ϗ�Zs�g o�̦>x@"���\U��d`�a寣����6"N�U�8�#�*P��x���'w�-�i#էҘ��G`��P��ymr�����G�c�c ���){��j��44����`Cj�w�L�oidX���4�>��_��]�ؐ	�s�e{[�ƾk���[�P�)i�!�4����1:!�f��).�o�d�5XH���bD?����R�O��X߸>Q���R2�6�;�a�Ԯ���.�E�u<S&�ӟ�n:�ȋ������|k{;��������ƀ�x��o�ÿ統���$k}���8�*}��w���ԧ��X4<���u�h9n�#t��f+�x���[�6�f��p�Fa�s �6}��+�%]���I1d�p�M��T����B��+�I���� EV��*#R��G�"���/3 ����$�å��*���y3�)f?��EŲޣS����ل�/u��٧�r��˅�2�P}]kAR�7�]$�Df�A��S�r^w��"�۪`b]�DEaI/�����uQ�A�5�ua=�D>\�VF-�u7� 	#بI�w�@7����"0�M�рI�������'�7̪B4=���՘g@�9Pۃ��X���5*�D�MO<M��c��	���[���ɦi(�w�z!�Z���2�?�s��cl��B� �'���))�Ƨ��gL��&�����C�ݗ��DB��Ƅ���PoG�?�7%l)("�q�F��A��	���S�g�ˑ��96��j��o���EH� �0?�a�{����5М�6�zv3����y�����J��qK1��D߈���w$e��U9�EQ<�O5VK����=�'�P3�/��7b�*-�����L�	o�~U���P�9d�#�R�q�0$kc`��'#+Fl�,�e�ܸ|P=��GU���i����q�CN�_7���LjPHH�R]$>A�C��+���7�e?��# s��]��J��h&�����#'솭�`q1�� % �l��."��i��M�F������:(�> ���ʊ��;S3-eA�fڍ���?!LN�+�s��T���1�qhf���̂$��C�.I����M�(�	J�b��`z�ƕ9U^�����w��f'͎�/�E��?C�'�#��G�[��r�h4�A�g�n�'�G��9&$�a#��Ò�m���l]�J���D���ƥ�������o+)���ύ�.�u��}t�p �ݸ������ۏ�t	_ p�eIX��l���ױ iE<�6UN�G1b�%�_�A��$e��D$�]�;�{e��[BS����+V�@�Ym7����w��K�%�[�Wf�%�;g7��+)++�\/�3��X�/�N5�~�I�Ӳ�I��??�r�B�(�GF9w?����BA�y�������p���Z�_�K~|O��P؅t��{�UC�u}��R�@������FIk��X7��,`�g�CA��,�f���

R��F��� N�����V:��mCH�2.�������/���B�?[�h��7�XXW{� �&wꗿׄ��'�!�V�b;��}GEmD*ŀ��&E������..?O����S+=��j�a��g��b	�����?(�u:� �I��|��=雮5����ժ{#���j�Y���b������i]�����b����uo��d�O	;xK&���h�p���֎J��w62I�Л���aA%�$<iȌh����'O�&[F"� �y8�ӡ�_�� %�p�dךM�^�O���a�Wv�����49�2B}��3��'QQ��首��|�Gs��2�sL�{(
���9G<�iF���Bi*
�����ԃ011�iV$�y_��w���
���W�n�"{O�6C颽�t��npGS��:�e��5l�����W���2r%i���28oVyJe�7nJ\��� V��P���[���K��ϡ����wv XQʈ80W5����khH2���E/X���Fyxss!��c���:��ܒ��mV���Y���{�}JIbF�S��������57�J��x4���s�LK�:��H�󕉒���c�v�H<��-R�������uy5�dʖ�����I`?N��|��$<�+&�G�.����"��I�%ƚ���o��kh$��W'>Q$[��{��������QY�xd٦C���J�k�o1mV��|뢭�dg�3���ԫx0�7W��Jf�iW�/(��+vC�Ba��G�� �GbɆ��v�׌S����a�ʋ;�:"~��^��m�b�䊄��{;�z6�5Q���:�{6a3F�p����d��f�"��nP��֫�:����7�a�&�pڒ	0��~�߀��ks�V:�Ne�zdc&�s�;�t��9����q4�h m1��ě������K�X'��[m:���O2�]sZw��W5��G ��?�y��H��IS�&i_�a�ۗU�q��)(�s����m����w��2+K���Q�-7<�,�I'�7��di.���+7�F��/\���q��Ôm�x��.�e
:��Iݷ��p�Ɩ"�/3k/Ȇ<o��9��@��4�о�t�PTv�:2�d�K�	�������+��#�K���'U{W-�Z��^)�ޗe5�<�@�����z��)���,������>��3˹r5�i�%�6cI����e�Y�5�$�#������I��^�lRb�K��� Q�R�����<cY��e. �F5L�.v$����V/&��4-�D����d�����s�����oRR�>Fh�5���s��/�ο�$�>^��ͣ��
��A���}Y��8��ݳN����4YGmN.�R��T�ύ�3�1��47M����麛,���� �&t�RŢ~g]���긇��To6MZWj��� ��K������=U���y�&���I�񾠪�)��Χ�'�� �O��d}����fK���5�)v�_�^���ທ�~ջI�?���b�g����eɷ/�y$-��	b�|�;�)��m<ۼř�-�,$�����U�^~n�8N!PTmFf�[h#�2�2��!�cx���o������ص[�²�;b �mm�#����u��h&�]��23Y��r�$]>�"�P
F�غ�Z��k�}K]4���Π�C�t���j:+�>������p/�3��K���*,.�;��x��1��e��i���
[X?��4�Y'od�����3�A�/ #��/��9��jT������J��*l��V']@�w��_5'ۺ�{���igy�J��b>զ̴���*�1�n��yV�l�/�^��E��-�BL���מ>l-p�ߵ��y����x��䖝��t�	�����>��"�����;�HOq�H>=�z����;|���%���C���3�5�a�{�A0n!4R�
�4���2��/�
Z�96?�~�M�[&���� ��]@���գ�ɾ=p�KD}T
�+��(��RZ3�d�y�^��HZ���rT޲-�\4���oX���Na�1�~��6"�JH-�L�C��'v&gph��rJǺ��ܰ][��q�B��x��]���J��.�����
ӝג׼_<�NшDq�OΞ�.��/R~_��f�$�gG�j���ezp�(v�pӕ�#�����S�҉����B��k�o�01��k�q8,M��e��cM�3�S�g��I�t�q��L�e�@�3�?>���[�c$��ӳ�}�_�(��s��-��P�(j���#׎*�~o��u��$7��4E|G�I���T�>�֮WI�%�O�hW/J(b �L�P�POjn�c��TQQ�n�YL�v�X�~y*~�<hS~�<��'�O�2�n8�7�3a%���F���yo�h��<#4�C�:�gM7�u�*}�������i�3іl������K�wݙ})��/oڽ1���{�!!!�n���
mXk��i����'7�윢���UD!�n��S��0r�Ǘ��)O]�X��S�V��SW�
�����֏N�m�N݁����xu��m'�DW@��5˲t�b�D��)���M$gЪ�O��0]�	|y���rY����w�����Q�P�dޓ�Kf��%��z���B��Hj_u�(6�?%+�����>��պ��(���c���c-!7_��"?@��4;���)h���n�����RG.��u����[�ځF��j�K�	n��sR斖W������f���`�3���qP��ۡYV1��k�E~�Ry@�<�7���m
s�����n@����'M�=�������M����:n@�R����$�t2G�%�������]����#�%��9ZF�J��k����C@ȡ���u�ۓV�W�惦7˾�C���=����O���ײ�C
�K-�.M�d �1^�"M�Th&o|�V�\�+[!��o� ��jUt����V�Z�ݏ�:��1i�YбPӥ�����3@�����I�W�����l���3b�3ɪg���xa�/�nu��M��[6�{��W'׭/
��ݞ����k��ϵqE7z�B�SI�f���hfP�jK#�՞x�+�b'��j��������6�yF�!���J���3�9��$���ySMr���,$cK�2��͆�;������5۽��wD5ka�Mя�5ǌʲ��������TbS��Q��1�io+��.�:��[_d;��`��}���^�^
�_-��8|��X�ӕ�Cٯ)�M���b�<���d42�r�
�~�:��ل�5��b=�V:On��"3��"8�:(���*
G�L�j/_�*��7k�X!�קP#5@�3����!�:ǃX��a��V��I���nI� �DK�^MJlcꯩr+C}�����0> �\�>��l��� ӷd+��c����^0��Ws�#��wH���b����M���Ss�jN��F}��	��mK���K�o`�B��7Y'qvv֕�-�t��ir�k�Z{�^q�1c	�۞.!)�����p���S�MqfO$�u-W�Te���{���LJ���C�}�����O��Us!�}�����֖;u�G
Tör��OD�Ћ��"��s������"1Q��[<����aGE�LZ�̓j�����?������O�'A<5�JK�;�_N�1�jL`�����5S�\Ȕ��?��7����M?~�|S�S1$��I~V�~��O��k�b�)���P&gF��qJ�IT&A��P�":~ąɷYI�a"m{�'���$�@����Y3�D��c&��tw$�p���(���S��4DS�Jr�r��D]��'�}H��R�O�V}dPL���N��9���@�o-0qi5YMgao�l��b�w��d�MV����Kb��A$^	��l��ajS������wC�� Ș|����<�	b��吜o�?tU�� ��"f�c���#��m�s䘃>$Sjg�5*�̘��ǣd�U�"9�R|&&2�O�lo���Ri���p�����?�?i��=Z��*L�_鐴uX������^��f�H���y`£_'h�}�f�����"^_T�92�wl,-��AE��N��&���
�#'��;	g�g�O�������~�/�$�3�z���zT\6(�F,J4E�n //�cM&>~��F���C�����p�O0SP�ɾ������	ǩ#��t��e0S����[ּĻ�>>�>�n�L�<Ǵ,Wr��	>���}[�P�'���j��5���=��Cl?ȧ�p9]�-T��ء���J�d%0���/siej2��X��M�DLu�:�����>�r���]�V�9���ߙ�_[�=���yɗd�c�����I�bA%�Z2':�~��<Z��Ɣ��	��B�s�t���F�Z��Ֆ��(��㮠�:{ZD�Sq��F��>��9ap�ᣉ;�|"�4����Ȝ�.���[V,dC��;أB������U�p��&�2���R��a��!�k�\��M�jX�'QN{�K�l5:_���-֒;5u�ᦍq���A�i�
�eH��H/}��3}�mDTCʡ��(^X�$n~�[=�A��9���>��e�]o4�&�O����vbY���&��"�7�槩��yRB����1�2������Ml�D��Q�e'����7�8�%ˉ+D_h�$0�F��U����bMr�qTz�s���hV���1n$�ꨣaU8�),�\P�aU�OB_���2�qY֗��ɯmVڟn��&��43�(&����}��x��c���Q S���
��y!�2��\ϷC1��N�wVѢ:�`�3e���da��i U'[�����[�ha�����N�N���'��x]H��S��W�w��L	:CG�	�H)�P�?9
:��<�� Zm?�Ne�����}uySzcs��5�d�ą#;lOf8oK�s���V������Y۱�����9b�ܰ��'#��]�%?�i�h>YM�k}��չ�~q�Ȉɑ�H���\L�D�7�0��C:���Fuw�4H�λcZ{�I�.�۫&MKE��j'I�ʰ�&U%*�9@���Ot�e�H��������1���}�Z���E`M��.=#
g�InH������U?�rr�.ħT�9��9 aq���N�*�2����A[2w1��R�q�JͿu]�T�����1��vٜ��Mc!z�6/��ʎ��Jq���W���"���Y�E�iV�F�̡$W�j�ۋL-{9Ǣ��ֈ�FS6��9�m
�:�9r��`Z3��Ywr��N�j1����%�r�����r��ӆ} /��D�9� 9"_�Q]_�:G���3 �p���Ϥcࠠ6� �OD����GޞG*��87p�^^)�lm�5��Q��-��fޣ�H_1
�Z.eY1�����P�v�oy��
���r�X�RN�}�>C,H�Ԧ�����E��4�x�|R��-������!��n��w�����f,6�A68��YSQ%%�d�|�UR����3��ԝRA\�|v�y���]WwJ�R'=+�(+_�̡.X#��2�:kɆ8���41O��q��b�a� � ,���0Uy	{���j�y���C�H �6ϠoɈg�Ą�}��R����� cL�ʀb��uu���w����SL�s���J&�4��J����w���"7�F�����]a��j�$(k,ƛ{sxM��p���B�?��C�H�GJ�ŋ�y�� �Q�I��>2�h��CWm@�^�`ڋ�t�x�t83�&2ڟ&�x�xTF$"'��+`e��a�����?��D��d�0½ċ��wê�c��n��nx�~��������'�ёZ�bZ��c#M�"�C�x�ˎ��~��0TA~���]Y}e]�)�Q����An�N�zyQ�e�MQ�T�`��<P>H}Y���\��e��k%�jѧ|4��*�g6��{4&ޓ�՞�
�fEl���7"]'1�2,���1�3V�:f�I��yh��h�i_�q�n7Ȃ����?���F�O��;�h����C���ub�������JȊ%
�LS(~/C6_'kk얞��>в.d����+{3����b8��qZYP������F��y�J���_;eޯ��-~�6�R�A�����^�{Yb���������ؾ#�i�W��M�r���o~!\k�u9ף�*�����iv�z��M*m��.��)��,���{��d���=�x�]���q;Xj�-=c�Aa�$���;�y�h��6�Tc*��G���?�u�1�R��x�s�v����?Цs;1�a�����_�2�\�'����B���;t���Z��	���	@$Hf��+�1���)����>��͖֋��>�]��]e�(B	�z�d�.a�C����7�-S��W�a����~��&���p����z�V� m$D���Ѐ�w��
�Li��MT=�p*�L�E�rj̹t���M���BM�����fK*�*�Ā�-��WX|c��"L�%��:��v���W�"��9�`��[��wO���M��_9%�Q8	PR1�5q[4V���އӘ,f�9�/�y������g��F�;4�)��ϳ��S������q��)6�^ØǮ/ʚ�*W�z����U��il?@8�^T&_B��<�S��$i#�O`�2R@BNH���Uk�N�*�+h�Υ_[I�9Ȏ�@w��O��X��U�o3��i{�������I���~�zqr�Qތ�8L+�K�Q���h�k�xȂz�g>�b�;�����-#��
�"��8��5ֆ�8׾��L\�(O���8�*�鉌��Ȧ|K�������(cZ����dv����Y;ˆ�."5(��� ���p��=�������,kՒ�����wr����"����@�grF�ێ�������}���Q$G�t.T������@�aɥ��|�%� MiՐ�k=N=]/�L����ӛ�&��=��%?'윳s3�e��6��>K�'B���f���|� 5_��躂���<��AaL�>+4����M��s��OA8��b�������!�@���R-\����0U� �B�I���T��2ʙ�w���r�)�����S~;}��q^K[�>�X��[ݷ��ωnV7�Y���~��D57��Z?��_�O2nʸ�x�ݞiq��-vk66�~�yn]s�x��U3��B��j�ˑL�C��.�φh���z���	�S�2�1�5b㙡�ⓣ�����y���8��� u���]��8��A���b��&+Ԓ`�D�
�-`کI�jkq������kF��1��%�^�G_�L��u�F����I�?P�.#[-�)�>�M�m���tc4���������(ZQ��#f%M���F���I�g䄲zιip�����&�b��u�ۆ�,"ߡ��+H�
�|,^*���2pb!D��i������^m��OF�`᧹b���!,s�v��M}��l�&V��fӮ�����Շ�yV{�PK�.z�w����M�5��!���0�JPu�@||\��s�.���`�~~�4`�kb�R8o)]�oPfss�:��p xӫ��G��%�Ҿ�2N6�n����ɳ�*�����
��}�$�yџ�ow3�ѹҡG-�ҝ���Ux7-��f����n��M�2�G�:�@�l�BGC��3��7��Or�e�t�4����Zľ��M�����NFhfiJ"�(�� f � z������XY�ƛ0��2��]��ؠ�G��h�-Y�U܍�IB���e�z�o�������*iSm�G��Tr�\�5�V<>}<���ӵ��#a�T��ڡ�����+���<��D��Dq\�J�{�
�a��4��0�P��q�6$h=����鬕<T0�KS ޭ��8�j��d����zϴ�WhW��;v�An*�8B�۴H#K�|y�e�6K�뿗��KW{=݃�۟�A99�е9�\6��+�6*��0M�-��k��D0���+J��>�!M�O;ש�ܪm6(�?7�{�i��F�{���!\��a�r� 4ŅX���Q�D��)ۖ�G�:H ��=�m��n�u �X��v�N�ǲR6����#�R��#M�e�vY��r�l]�L�D�Lʒ 2L�*l��ɘ�HdU0�u0����M:�[�����rY?�
�a�X������F���|��j��n�~�R��Pȫ�`�VȁT�2�0JT{����2�:�i>=�=����r�U���0�R��
�CrƗv(d�΍& kƭ���*��|X���f�ۙPiT��ܩ��� +x�j�y� 6��eM� ��N^S�����SXo�eL1�0���Ay1�*we$\�
�^	��Ûw�u�řY:�:�4t�-4a�	�O!HJ�C��-��]�A�B>	��Mq��x&��q��"��"�0	$D�(i�4
�l�֧�Q���#j������~|yd�{w(�%�{� �{�/��<�'.O<�AK�l�>�>�/K�컼��%�G�b���Y�OӍ���{)�`ne)N��,m�����W�)�O���u� ��)'�,�`����pW�'��q,>}ADJ���![|�ŉ*����q/�y&�}A���o�j��25�Q�3��ٷ}=�q_�Q+\���g5:l��}�+fM1��4֓!m1�bQT['�qڶ�#D�����=�<dɪ���O'׽��'L!`7�)�;y��N�1Y'����C��!��֯�߅�jq�	z��E���H��YX�Ym�g����	Yo��Ш�*���X!��)����IrWq� @�f_nV.�\l-J��*�
�$��B`���u������FeQ��C��J~ǾL4�������
O���zv�2�q�@����_�x��\.6�������E����dР��=�2���Κ�c�7?��&D�H�f�ؠ��F���������h�� �J���DֻZ�Y���⹇���<|�OҪ/�ab��>�gE�f��R"Ỹ)pҪ8�({2M��WOG��Lc���B�b�:U�r� �}w��W��HM���	�@���>�-��lBvf���ڵ��W�$$��qn��ٮ���5,�]l��� �a�y��C���
~\�'/~�Kx��JSZq����8yH���)D���H��,��(�#y�W�!pwoɖ��Ʒ�:d	�iR���DJJJQ]�t���w׳��V>�_��'�X��J��F�s�l�m���T�<�g��v��סHȓ{~�8�:�6r0wewTأ�w_��a`DY'i�V0v����$ؗ�%*�9�4;&,�\��"C��@��.f71�;C�# ��[-�p����.`�`�j�q�jܷ�s���0=������.ځCu�)di�2QR��HQ��]z�6�wFJ-|̋��<�p27#>��Z>�4����������ml�����O��h6�����P��pۻ�o�Qc"�����Ѐ������y�or�7_a"vd�u������,3j�?���;T�7pSIҀf'b��\�Nr����6(b�_����2h���L�O6��D��ǿ��>���k,�\)9d$[����u�$�%���*��RA���?��:2o�ݔ��Vk�r��A���ʿ�(���L�J�Z#r�vv̽�������w5��"y?$�p�U�c?�!.�5cl~�S�p���c�!������_�~)G�w�ŋ��a����A�&����sBh�p
���>��<͂��ݠؐP�4�N���Ç;�̣h�
$^�ȕJ,����N�ٵ;1hjǤ�ʰ4W�����=�'�#�㮁��.iyB�B�%@��.u�&L+�A�=�Va9*md�Ϫ�Q�/����Q�]���YCM&x�P�^4��3�El�k;huȡ��3�A�c�;�`��R�)�y_�:����t��\V�G�jW��M���Ò
%5A��G��q�g��jH_������`ggf&&���GYN�d���t:2�ʵJ��I�?���nٰ��z�ogC�a����P���_���.���h)��=L�����bUP���߶����l���������>�OR�!7z����=���/�'��p,���m �͟��3�[t��X\�|5W�ݘ@Wu�����D�c7�^s3[N.KEuY��>-1%("���M\
w�6��=s�o�'�{�tH�Q���-8�%n���ℿ�c�x}8�LŦ]�SGk:J#��謪��N<�����z5��]�S�y9�`��t���<��Ĉ����zO�8����8�{.s�)�@pS�ut��1	R����"d"#�Az�S������(�4Q$@�l��N=���n[ɤA����v#�ᨬa*��q/���؄7���@����DKuvU���̟l���<�gk-*�pݏ��2�yp�=��m��\�t��r4g�[_���[k�8B��r�&g��.�f�c���.x�W�u^'u�Sd�9ڲ�ؼ�Cu��� l���*���%"�s�F3�w�ber�^n�9���3�f �y�-�'�ޏf"+k�9�S�����Sf��N�>__����e�L�+�Mpl��9�Ѳݵ�3�5��=�*x#���Y�QG���]r��k��!W�3b�?�'� T�kF��Yg��׈���Ѻ���M����ٰ�k���Ѽl�z�l�^�&W\�~�N��k���ҳ>��`��:��`�\�V�}�k[ܺx��3� p^+8z�4j9Xs��F�%u���(�[�;��DȄ�OM�l�������<*6_Plv�F�D
kSz^/hW诬\p4��qXF�����359��UH�,������6�[�/�K�_��<��5�9���oV��tBM7���Z����w]ޟ������@������J�q��,��i/���z^�"��?"��rw2?Q[�u�%�2�כG:���O������J�}<��]ۙgdy�.����ͺ7o�m�ô4kѵ���کe�~D�������#�I�V����Е!�f;���Ɵ�/[�t1$ׅ���e��D�v<��y���O�i�ic�d�o�:����8��&���t��_����X�0�T��^��x��^qu1L7��pZ2䂗~�!����DbBmʏ��Ʌg06u��n8�۲\��iV�ד{�9��(;pg�����r���c:O8W�ƾ�"D��stu̿	2Y���d_�=s�_ӄ��,��S���p��I+�l�!a�<k�X�X~�$h�ƻ!�	A,�d*�Qㆅ��x��6��£�Mm��o��s�SC�x���p��6a����b���)�$[3ҥZ�a]EŅ�5ȋ*�.��cҹ�Q���ި.��}��@ҵ�8c�~�5!�d�1���T���y��C�*��/*�v걝�*~��:I����J���ѹ��ҙ<dg?rڱѰ���B"����f�A�-���xa�/v�X��ưf�0�v��.����f�N�[��g�W����Pz'�h۬�����O��*4��&���gtӚ�X������ON5{��g��v7��9�	p~���t!},k�������9e���N���Qϖ�����>�|y����|hzGÉt*G�c���9�Cq���U�z��l�g�q��h��$$%�F1q$l{QT@;�6e�l?s#8B��=�9���0����X�	���VU�j��g�eN��k,�$��qD�$zmW�t�Ӧ��`��,�8�m��7�_�@��պ���5 韉�n���Β^wK�ڛ5w����@ܜWo��}]c�j��;��D�Ӓ��O������u/�p��1Lr� ;'�:����%��~LD����D��ܟ��b��`�5�,������8l����Z�4d
�oLen���י�xB�?>=�RM(���Z�ü(�z�?�|�Zּ�sZ#Q���h
�o�2�;m�
['h�=(䔞}�,N0��~Rj��8%T]Ag쩑x���pO��SK�8<��l,����gT�&_Kf�O�� I/��%v/��F�����c���G6��Iڎ�i|3���)��j�E�`�#�[&j�0>�37ӌ����CV�H�=P�X#�OT|��
V	m����?��>*"KV�s����_,Q�VTx���|����\����[�;�"1'�m����i���= ���*�x%Ґ�m�
�����M�����SQy��U��歉H�7��yr<�1�&��Eg�naIP-:-4��rRKU����.�zT���`@U�2h�������ة�%�eg>�K�E($(�f��j��]b�٤�n�Eh��U���x�Wa��1�C}����<W��!��~߿承p��Q�v�����d-6Tks?b���I��
G=��@f��#ې��R�Y�͢�ɾ|���P��9�u��GD=v��q`#��%u�Q$�^�ir\�+��F����{��ь-T��Z��3`	4\Ǹ.�R���Y�|hд]�h��ct�Tw�<���k9+��`�v�zl��ǻ���Ӗ��GԆ�n�cF���߆���U=��5|�}����~�jL}�<�vf�h��s+���Z��;EU�^7a���7�Q�[�s���ge0��%�a����߃���pv�z�5�n�����1$'0����s�ƶ���Ⰿ)U���Z����f1Q��m ���?d
*^�|����D+��Mm�wYj�b���wb�{_/>�v0,�jPq�Q���? g@��N��qG#W]N�������uLt���`�7B�q����?���r�K�>���`ݗ:��}��2� ��C�)s3Mʇ�X��h��D7\��Y"E�k�5O�R�]w59���9Jv�z�};_�qS�e��o'���t��{�غ��/�]�G�['�S/��ʞ�>O�_�s�:7�x�-���l�~����"R��J��д](�d1��/ ���tف����ڍ$ֺ�Z�?7]H��ڟ_eE,.%g�|��>Z���'RN&�_����$ρ�j>�^�?�E^׽H���sa�����������G��g$9=zF-���{�c�h�}��29�&��?�q��Sӛ�xʣ������Y�5�+�����Fi�܉@�,њ�)�*�p�����-������u�������uD�t��UA��s����l�)[����~~)�'}�h��YT��z��}��#A��}쇎ph׉�ɓ��Z�����%Y�k%��@��vqhdA�Y���5R��!>�xQ�-�M�0y>+��a'�*�F�&���)W8��DF����<l!c8>�]9f�4���!ǯ���=�4��m�e��V6�n���ѰvS����_��-cAc!Ģ�����1c����s���d,�8���ύ�1��ӧ�%�vY��ïy���|�W�5��a���}T��Tĸ!�Տ�2G��]c���9���	�'3�-�,�����s�z�2�1�l�%�sf�G����?��Xd�@-4O��t�@��тnp�a4�7F4��)s�䇒�?蠮�����]�A�䵵�$�y��	�A�un07n�Ƒ��cH|���L�P)Njd�[�;���*���O�2��\�'�SO�niƊ�¬��n�gi	����h��_����F>�$���L�+�ܛ��"5g���3��(�I?8�h���ߎ�Wu';�89{-���3�8G.)t�7��|��$���f7J=����+I93�U�H���
�?-Y�9B���^D��F�[
�޲�9\�:�^R�Bt��D{}#������Z����4����5}�y����~���p�I�^�%���r�;LTe�~��N�4���uk}O�.�� 9Rt���s�Fp��Sߏ3~�>ƵWQd��0H���W,�9SVߨHU��)�6�}����~~ri#�&��(���u]2S�??ҡ������=#����ې�����qA�y�uy�?�޲��j�Z���{8�"�w������d�'�G��/U�r�J��}�c�˟|�����9Q�E�U�����2���}s�Nt˜� �G��z�-k�~��H���@a����#��0�'��H���X�8["�%� a8��-�f&c!����zJY�#r���oy1a\���E��+�d�xa�J�v�@3�[���_e�㬇�`�Ǉ1�܃]'��`�Z����*�%�Ks�8���Nڑ�_e��0�}����j�[���F����vl�4.��R���Еl����E$.4�F�`�0(ccR��C־�������j"cv#���I�с��p����"1z<�ˮ���þz�&-TC������u9[ݘ�kI�C�>ң�b����/,'�J�NW���C�����l�*/�(��z}�pr��7z,9�v�e����'Hq�F����2#��u�-^xN
����R>�:T�7e�k��w�^���{b��몧D&�r~C��Ա�G�i��ƌ�5�G��B�T�/q�U����O$z���$ŜxS�3�G�SYAb����ˊe��cI��Z���]x��V35�ݛ��k��D����,Љa�x?:���ǉ�ja������wig�z�5��^�|ɺ���t�#�N;�B��N��D��Ia��-�������v��k'�j��0A��f��?<X�wL�C�C�7�G�Ӄu���VA������ġy�9U�=�@r��w�Mw��U������l��:@�b�m�'��\#}����"���)n�������&A��p��]�hh�|��[_"��]6��CWΖ糃C;����d3���es�&��8��HvEZ�pOoK�]�0h� /�D"8"#���E���-[��'��Y�lL�e,O;��r�-�;!���c�)�3�haL용��׮g��ǅq�C�t�,�81�����{����ۂ�>N�a0����ec��4���z�ͮ��<UTTP2؊6�@e���st%�*����ܕu� �|,L|��zl��~����ج�NQ	��5��vJ,и��?P>��ͪ��Q��I 1n{�4誯(���uՉCH���w�$�һ���@[�(z��!{S�^�nl#���eWPh�N����B��D�-wУ�b�Z����Z���|�G���;�
���\A�,^�~�t,����?"1ehl/�����w�����&���Z��|pc�z�wښ��(�~��z�9�}����T��n��R��%|��?� �s��1�-���7&�+|�T����5��:��9iK������ �o��_��1���f���]F���L�A�B>���?���F�z|�|_?lv�?�P��{�r�YN�gz�V�i'�P�Aj�~���~��#�w�Aw���F�At�3D/���O�N��:g/��^x�Q�r�.7,�ڡ���:n욚P������}s�ۡy��G�� v���_�Kq�GA=��e����q#ѵ{��Jo��
�^/A��FI��B�Yl]a�e�d�ĉ;V�\�h�v�~���}0F���Uf@���O�o��-��[�ٟ�1�`��8�ޗy͂�Nf[�9{s$ZYm1t��s�Ϲ�%�����|.A�l���m�3 ]E��T�,e��d�&       (Lr&�~*�1gN��c�n�]D�3r脣�>:-��>�Y�,W5Z�ۓ��}�L/�u��_�ME�������h�{9�����D�]{L'�F�h�����y�rv�H��Q��؉$�Dt�H��V5g�fr귒s��$��~�-�$�z�z]���$xt�-HO�`�ʋ�9+j-����'>�������~}ʉ<�G�#O�u>W�(q|[?+��5L"u��m��U�CU��Q��|aw�s��7������5$Y�^;���&s�3ORh� �����&C�$���G�������i��o1\���W���ʪ�Lٍ���v�?'��H�jY2�/#:h�����Se�6U�]*CS��6��n���[cS��.$��;ߵ�&b>��4~`4�,{��Q4��4yK��?�W����w��p��U�84ބ�p��Z�FG�\����q��f��^oW+w��V���ı{��5��/+��5th�&��l��T;��8���w��]�F%�z�߳� m�c8W�6�MEk����Ƕ|ى-Y��2T%��M�6�Xdl+[���f,b�2Ȳ�(<�;����ֱ�?�߂f��>�D�l�� Z��`��'A�u�s��1[�Rea��Jt��AW���ob�r�X����^B���hn��7ݸ�5�m���7�|"��o�3s?�>5R̜���qi�W�XN��:��y�5�u�H|�3E9�R������_)EQ��]����Rp�D�7W�~�����+e�!��+rֻ1Q�=u<�6��W~{�����ve��-#g�o�6g�r��66ES�i���&�0H᪲$nr���59m�:歾!z��ҝ I�����_�8�g3q��X�B3s.C��A�j-z�r7X�Mk�|��h��g���o��Ntǟ���$/��퉶Z�üע���/�p��Ns�U"mNn�������ֵ�ߡ+�eC���j&j��jYg�i,4g�����H�&�w�=*��$�GE���7���jA�o��5n�`�ܺE��)/���b����mvǙ ��(���c_�wh�j���$z������DK��6��0���ϱ�Y0p�'����3:1a��FtWE[��������1�I��^菋3�l�o"XȚ�:gsnv�9o����b-F�2�K�-�8��\A������3 ]E��u���P�`��$/�#�xY%&��\�p���"����dE��O��ݝ�ٜ�.��d��AAPQT��@EDEf}�O�,�Y�gBA�H�( iI�����;;����Wչ]}�v����9?���7ߺ���S����"��]I͘�;��դ|��MH���Sf+̻���?��o�����X7�R�[����I��╤|9�-N�i�Xx�j~q��l�	��a�蓎u�0_FW����6��!m��Y�~�g�:t?���[��R�Spt~�M�]�?_�]�mϜ���� ��˫h�Cd����)�����c��Ar�������~	�7{Vs��������swa����u4���4�v�9WK���xfی�ˤ���h�%�qc�i�è�U;�h^S�2t��c����l���������c��z���*G�+�+�7�s �ҍ����e�oF�m0v��r�;�h���6�i�X��)c���O�������^kD�ZM3��oeZDZ��blٲ���H�t�l:�_B�q�
	N
�I;B�Q���y9Sb<�H��}�G���3����V�֭���޲$Q�ˆ}�B��:��@x���]zl�x�@hb
CAA�6�$��3f�:�j�jo
����;ø������B��K�L���<��?�&=�% Q+�녳£+k�_w+i�G�Ft©n=�f�Z����H�y�=m��w�4<;x��<{"�aMen=F�)p�-Y֮��cL�k�X
^$���'�hn��h#�Ԩ���#���-��:��PRׄ-3�����:���!뉋�*�p��Y�=�ͼ�̓H��c�R� u~�i�.��淶��CJ{�H��c�z/�z� v��2+��=�\���K4<�ȫ����f#����
�	o��>�;�]RD��o���woG�Nv ��ъ��t?g�3뙪4�3�}�8�����;]=}լSіl����x�<M��,�Еm�-Ӊ|nz����^3��M�>붅��Mt�yt̘趷d��ǙDf_�t��t�V��~�h��-Ǜ}�(a�u�ِ̙y������f�����ɓ�\�b��oQh+`�6쉺��mJ}2�������_o�/Y��?<;ll�ŋݻz���+Wf�H� �	C ��?�i[&� ����ah������Oȶ��148��c�s��O�ߟ�3z����%��ۄ8F����~������K�.�9���a��-{�
&� �qvI	��ל������~�[H��\��H���c]&@7�p�52�1^0���F�]sэwEs��}�H]x�+�2�z��k܋�ԥ�GK�,�������Ha</l����[N����{�y�w͛�Xf]>Db�c�5�ĥ��W��蘃I���{��d�S�pX��iI3�
��ȍ4,N�3��)n��p�IS(s�uQfK��y�/x���y�HM�a�e�u��n����O���974/��{�^��+��S�>�iJ|��޲��y���d�zpn�IQ�:��uֱ�O�c�NSC�}uۓ��J����ԝ���wf��Se�@@�㦗���Q���Stum�m�Q��E�ң�5��+5��q�8� � z��s>K�e>����hYڇT����֚;�m�ݻLѽO�߽�#S�?{����l�3��������a{N�pM�}�8��^g�q�����}Ϧ��Xa읁�=/�=�"�8e�@��q��G>�z�l�{)X�t�������+������/D��MU.t����U�z�~�A�� �B��]�����̎� X��|��>�F9 qz����{:���id�d�n�x���0=����=r��-��Ϳ�n��O�[���`�_,���{�0��O�S;���9A
�-Њ>=pj+�~-�$�l��{��ٻ"/4�� �Ǐ�r�k�������h����ǾC��:���ͼ���ט�6#�p_��Xl��R�Oԙm��k�䚷�e?&��GH�ȼ	|���G�4��߲���/�:�mN��g�6إDw>Lz���_~����ܺ���VJI~��z��s"C���ޙ�p����\�a�\��'~�H\DG	A�,7�D����e�u���C���/�4�����ߏ����v���o�ü�w+z�|Λ�i�'�Jt��H�.����E�g����/B`n����系ڛ�Z7�b�N����Sٺ�� �����8d2ꀱ_�!�����j$�\���7SM�~օ�*O2����pH�[����|wEo8�m��ѭ�ާ�� ��c�E���!b`�f��Et��n����^�{;{4�6���fm�fֳ�M�߮�f�O�M�G��iǋ�Y��+��P��3$m�u�~hW]u��-�_k��G����1�g��0@_6x�x�0���8C��5�\�w0��IY�ʎ8�[v�QG�	M�(9��3��_���~��h� ���a@�?����~�K_����<�5�Ӿ��k=U��a��]�}�`� ����|w�q�yA"���袋��_�:��]����PIv����.��B;��#��r�kh��
����]�0x� �gKI��0���$Q���E�ꤓI�
?�rFb����������M��?[���8R�s��=D��H���]v!̓+?����C�@���;?�,�#�um�n��y����|�8��ӬO�ǵ*�	��:�����-��8[l��_��v�ÅIq�[��o#��RRmƊ����w�o���I�o���vx։u�)м_����1����f�q�;��3m�}�)n/�i3��<4
����4yAGv����������<8��3i������ǃa�n����_�z͉��qa5��/D^V����2�Xf,���"��<6��A�'8�ac��ݳ�&zˡ�UN�~�d��6���i��F����Tg*��lE{�Q������yYD�˔��Y��y4��Wj��L#�^I�]م�ikV��y��3'W5����vE��j�R3�~[5uv+��Us̓h�dM�N$Z�cc�w���6��?��u*J\��TW�3"`��s�=�z�8\}���������w�A��կr�����|�>��OZ�k^�5!z6l�@��������-���K�p�p^��W�{��!<BOD�����>��c��>�6�G�_��W$L ���L�@����\p�v�a��C!Dާ>��(᝼��O�T<������mo�������N�����=�t-+O<�^r	���O�*�#�����[��Yg�y��>�l����o���уG����źJ�~)��b�ظgE�>�������]�;��f�䰧�W��Uks�4�d��7�7m!��y�?q/���I��p�������[���i��[�s��H���� R'��w{����[�v�>R���]t1�qf9p/#�5�s�5te_�$�ƚ�8��'W�ua��w�׈��n�%�v϶j�y��H=� �K�ˇ1��t�=���s��l^���OM�4����bg[�tu��ri��5� �goٖ5�ZB���O�5?���t�\N;=�x��s�(����ڷ]h�f��gW�v��8���@�����0�������-#�X/#�Of����a���k��;-ރ�տs˭_f�㤜d&��g�_`h�:~j�����1���A�k1��Y�5�X��ru�3'k�wEs��;%ܜ��F�]�{��v7��Q�&�ޮ��7��5�������f�Wg���?����<���>�9�)��m�,��9ìcb��3��{,�#0�h���Ӣ��/��W�a=��q��/�-�~�鶟�PbA���S\��!x� �XH���	@ 8�裏�_��6��P��lK@��;>C��b�r衇ڰB a��������u�K�{�WZ��e��>p�.LC<��ڇ������7�t�{�w��=n���0�>�_��e����=��;餓�4����-����%���m.|?��l��K.�ĖA�Cw����i��>��E���P �A�B_*�A+�i9�-��+]������~@�t���=b�b�2�6��'�8h�<3��c�o�I$�~����]�	G�ڲ!w�)��~��ȶ�}�̧�0��:w��v3u����O2n�L�o�\n���r���B?��M��8��;�!��?�<'�J4m*)H楧7�}��f��}�m�н]z��k�>��>�y�o���Z�0&Ēw̿������G�hq��4g�#lA駞r�`_w� �����ٹ�&�PY���D�����f����؟��V.7�ڭ߂�J\�y����>7��>���Z2��&�����,wIW�.u��Cq-w� �l��:�j�Z�x4������c2˚s����Mo=���]"�mA���>ͅ���f��`����D'v�Sw����I���湗�n7��fm��z�<{���`p�;;��FQ�w��|��'^�Q�k�)ʖ�nq�HS���?k��k�s��?��M����o6�y��yd�[��Е�T�9c�</�*jU�^B���M��nF[��پ��F�YC�vo�6�>�[�3z�y�u��uǡ��-s��F赸��=�p�3�����i�3
��T�Y�P���0Q�1?����殻\�j��G $%�	ĬY��s���򕯤�ow��<�lGyd��}���X�p��A99�����_�9���s�=Qh&��A�k�;^�g�l�hD�"���O�i��ñ�<��,����\'�x"=��{�b;���?����K$���^5>�xH"�j�I�ĺ�^�@ ��5�jC�}&$0 �
-��UF����]b�]s�|�>��D�
��2{���l��� ��\R~�*�*5��F� �s�~Ƙ�q<����d��}�0��Mg�n��Z[#�\aP�K�K�?�tc{)�t��`�9҉@�'�e�"G}�y�����a�'cq�|Q�t�a�&�~]
i��t�,�x~ڭ���^�������`�x�l�yi�ċ�O|���P��|(���A���~�E3�� ��w�V���ߜ{�2��4�����f��U�����4i�w[HM�K��cp���<�n1�L/����O<�ԦuN�s6�C#`�~��kn��e��������TԘv��7Y���z!��˖����� zCm~(����~�����N�Z$S�}��mޅn'p87��u���H5���Mъ���}���;]p5e�Zl�� �����m�������M�1�j�po5���:�?_��#�}�f>�wc��o�6�d�A_��}ɯۈ�&s�}��w�6w�/�?v�#%�V3�߆�͹X6�^� !�T�a!���O�nC�84��S��%�Ʌ6�A� ց ����za���P(+�O�Eσ�g;<�s�y "�geҶx��{!���	7p��.�Ii��3z�,���D�"���Kʢ?x,��@@b\8�.���n�w�0؃����X�P�i��e긅A��2D�*�3�@�Ʀ�O��nh#2�gI��И޾��F7�
���\�F�`�(4���uv�4�ÎSf����kh�`^,�:H�q����lYo��UT�u!U�I.>��I�|�!͚A���H��ٯ-�C9��5D�C�	��@X�8s��� �^������\���%��5��� K�]�y�p?1�;�ц9Fi�{�\f/���J�s9�3'��|)�\�����Ƙk�D��Ny��Ȩ���6��A
IS8]������������yiS76��3;Xg��	6���b��v�Vg����;��Vs]�{�)�=Gg v��P�ܢ����6��p��JnA9���FR�֎`ܳ�6���:-���F���m��������T��^mN����^���fwj:�f3}���NR���>����v3ӯ�ۭs�aw��j����aSm�����4sK��-3������v5��nn���~.�ƑZ��Ӽ�-U�;[�خ,�������;��d�ɂ$��%�
�����V>��b��51�5�����rgx�I���)�����O�2�����ܻB2e��a�P�EY����^���U�pW���`0�i{X���֐ �0Ʒ���\���9ġ�[�F��M֐߰&�Ol���O�O?�a�9�81�{��K%<�p�|,�-�:&��{��}�Y^�@��;��O�y��4b:��f��W���3_����A<!4�@�	O�	�BvC�[�t�<mސ�':/�=�k�{i���AxC��Zۡ�n[�.	Àd; �C�����b���"����*�i��� �
ƭqHg?���O+����s���Ҋ^w0�k}�;�V��l���3�7���r�����ܘn�=7!X�%�����|�F�x���	H�k���L��'����S)��l'�-*g;a2���W%�9ܯp���F��g^��9�7��@��6�)�gBrZyc6%Џ��{�bk,±��N��� ��0��1��8/�V����5b h֖�b��n�{X��%~��'�`:��,�����hȞb#D��S��$�pQ��s����ϛa�7�2�����y��o3:o�{�{�)�2΋�o����T���ή#�~ٗ\v��yP�x�t1"1���Adk?�VhŢ"A$�2}KZ�j3_k��������zM��l��f�PƔ�q�6M�}P���&��n�}�w��Ѓ�mD�*# ��{M��y(���;! �9��"���t���{-W��zJ�R��km��#�*�b�AZ*��d�nU���	.�֦u��|���Ȱ�W�d�ɱֆa����@��}�r��-u=��g5��hXO!�Ŝ/[6Fj?4���2�ҧ������h�����G�T���̗	���٬��@��6D���y-.��nNtm���ޗ�BW�~T+6|��!2���v����/�!��[gg'��6Ge2 ���h�w6�*��J�]Sn��|$&̠�b��m�Q�%W��$!vBZW�T	�J�b�z�r�+QO��mF�w���s
�����5ݳ1�M����~6��'�N�U��N���a AGs��޺u��3��H��j�uq�x���@$VQJ�\�ԃ&��-w���A(�x�����'���)m�>V�G�u�~l�ڔ�����8lr��D��j�
��#p����K�Ȩ��`�h\��2�⋫i��NjkC�0��v��M[h��.��h��M��;�c�,$��1߼eQgz%ߋS��[�*�f_�`�-����Ζ�H#|�n���aK��
OQ&q�ttl��"���?�u:\�j-�^����2�Þ��#n��X�"����
�Q�:($�h�C���K.�)
��ܣ��A�p�!�IB\T_�k��k��/�w_���%�z�4�&�:�j�+����ӦM�^XI&��D�&��&/���6m�L�v_�}^g4�T?!��l�8�s���8�&�#���}oXW|�4�_�mdW��)?]��9�P���S���	;��6�g3g�#A���Lse��X>F-h���b����T��R�iZ�G�\m��KƾV��$�)��^���@+j8y򔉴e�Vz��gi����ec�F礴OHY��ڶ>ӳ��+ڸ�����3�h���4vl{T�H����A�l��/� Ki,��.��1I��IF�"-3?U�9������ӗih���i���3�[��R$w� ��>0ƗnsMe���FZ߳Bp�T����<Am97�B�ߋ-�q�`S��b3GRð1^���fѿ�]F�>��-[�h����$��O�A �f�GՐ��V�ZK�<��}���4c�4�_BI4��zKm���]�g�R�3(n��\�G߼@mm�ޅ����I�}�����A ?�2���ٔios?a0�T�V�z0J3��hNd���j���Əv��1�sg����QZ��˾�M�k�'�n��5�oㄪ���ǄpGdu�u�<z~�
[��cOѴ�S��F���� �[���+^�uk7��i����Y�$��P2�j�IR�T�J�#K&-��)�TUP�K�ђ�_���@�y2F�u-ڃFa զ&�]�Aow4ݽ�BJ����Mgj�������;��.�ۛV4��	��'�Нk���j���h��}��!�zh��^#8\�T�c��?�Ikjj�]�ϱe��o�U/���k�����6��h�Q�F��H�_�!/l��������e�Vڶm�-kii�]Υ�����_���,���VלJ[�[!S#O�|�,�'��*{�@F����c�Pj��i��[�`�fR[ֹ�9��s�bS���bB�7��Q�d�ւa�����4��G&��QMn�go#zru��v�[��Ն��	i.�|�����Q���q�4��)��}��*�l҆)S&�4��6����Gm���ۛ�L&ۇ5g��	�YjTO����r�5��[o�v�b���q�e�m�ۯB�Th�r�W��_���E�jnn����;w�-��n���m;-	i�ҩ
��3�����$� � �P_T�@#Y�|�3S�ޤba�I޳�8J��k�,�z�h��f���G�ڲ����aĒ��랳�ݧ�C�v�����R�'Kiɬ�����T㬤R�z3��t���o}u7�r$T)[Ҋ�Ǻ��n7>a��=	�N���d泹���Lu}�&M�H==�6RBфR�=����h37����w#)1�P9M������D'��36&u��������]�a�B3��h�q�Ө˜@�)�зƇ]�Qq�u�>�;�Q�m�-�b�tG5w�t�c+�$��8c
5 ��˘?�ݽ�}�ޱ�V���	��C��U)�!ɦ5��$��[l���=ԛn�i���Zl|�{��LKKs�E�E�勴K��+���+MX�z�����'E�r����?����m�P$e�2�[��o:�{Pr�	�a=h�Xn��<��2J����� �1է�Y̠�IP�H��um�䋶�㣗P�cImX��A�w-�A�'��5��թg����m�w?j�6���J����_�O��Ғ�u���D�gWB��cm�S�M�.k�eSZ5���s�j�rR��U;>��N���������̗�Q�QX��HR��P-K�c�`�
�k��N3k�|c��4�yЌ!�b��L_u�-ky�)j���9�7��5>[� �/�����-���'���ZZ���-�H�t���N��0���Sj⡤y���۫h�(E����0Ֆ���H�Z� Hg��C<gg��@��{�EhMӧ�ZK�Ƹ����&jl�(�� ��P>2�i�E����h�j��+Ժ����!�Q�wo��&زu�<��l^G�w��Ng�=����.�1%/U�1u[7��sz����hZ��w���]���-+���?!a�J!!ǟ�3�g�khHSWo-��MW�2b�v�dZ��@�ZݺV���"Ԇg��8[��O����W��ݧva�^���=�J.� BM2$-4
�=���Le�����~�6���l'�\�8C^l��v�.ݳfѪ�>NS�O�ӭ����1�=� ֙�W�~jB�������ez�n��Nv��FZ}���g�|j�IATC��8'y��հW�Xҡ��!q�<�)Q�B�������mٵ'��}�L��k�ka���f�M�X1x\�$ƚ1�߲�f�q���c��As:)��&PyO�Xc�!'�PU�-�]���/�%QUb4�%�㍗�������2�׎唲}�@�j�3��K��N�_�;u\�%R[7��׭�������G��K�=�@mh`a��ׁ��<�@�]
}k�J�v	?�S��n%������N<�2'Zq�|�^(��2<h���`����B�!�(DG�vm�3�i���q�^���ߝ��~��K���'ڰe+�|֊��7'����PFy$��{P�h��6�;�b�m4��ﶃ�u�Z[���Jg��������E��JD� B�P}�,y:�Q�"�<�"Z\|�-�Ō'&1�1�m���i��L[��\{��m�h��7��]g�R�G���y٨�rr���H+U�jy�	d����&}���C��eQ��]��_G���|�b[���Җc^a�������YҽN��a�U����*�'-���yJ����8�Z&��ҙf���K9z��>~A]��X�ŊV���/>�G�
P9K�V�:��|�WS���Է����y;�u{l���l��Fw�{�8KY�gn�|���q� uI�ȃ	�R�g0�}�����CB�Z��N}�Uڽ̛�2]�p]5g.5�p�-�l�>�5�\n��n�	rc��"hy�}	�Se�|����[F7:k?=v,�L�J;�N;v�g�z��$��D�#a����{��+�
=�jш-���Ľ�,j���P:mD�_��y[i��[�mZ��UclٿV7ӊ�M��ӝ��w�+������e=�����Ǣ�B�s��m����<��:�[G����czh��ݴ�vz��.Ӭ�ǈ��Ί����%5B������^A��z6̫�H�Y�T�y^��X�)��@����XJ(g>C*nP5`�ϣ�IP��v�w�,�X��  ��IDAT[�y�l�x����͔q��{�i&Z�J�a� �������Xy�����RM�Q�XC:M�t6���Qq��,�U�G!���)�)� $_y�}]����à�Y�McJӢ)=���H�^E�h)�>��Gޗ�[��dQ��(�[��
�%/��wc���F���wo����,�r�wR��~�!'BT�ӓ� Ѝf���B6�Q�|$��R����&Z��j�-�T��/Ĥ��p�Р�'[ɠ�D�9�9¹�)�3I�G��5�ԢF�%��R��I늗���Sn~^W��K!~�֕�͗�[��0��;�cI�-U`:i���?~E}�[�}p�k��8��`9�ۓ��]�h9�$$���a�{��S,���Wx�|�� �_Jg�~2~�ՆT�j��Lʍ��2���1���]�=��O1|�넲R֧
��WG�-K���7Obt���Oj�ȭ����=$�H�o/����g�� Bat��}b�g���r�us;~j1B#�h�z)d��%�죒޴h�[м�(�=�quQ�5�PHc���h<O��#�6[W�>k=ik@Db������B�j��[��o�ʊ-W�(I�>�%i_��w9�Z�������J9ϥ^�|�o���o@���|d���ޱ��7I������Ҁ�q��-|�JD
T~�$=W�wޛi|ɮ".Z&�ЂK�1:������hWe��J���r��Lj`����s������PR�R����QA`\R#/Ң�To{kװ��]���o�Lu�ʀIH�.�m-�J�x��K�v�_���J�٧�BK.U=�
�B�G!`�Z��p]\��#�GPג�*� y�Z�>b�� >���M)Fj�ݭ��J�Ľ�Iϛ�����IϘ�gR����ȉ��W����夲|}��[&B��C;���$aWNRhB?�k�qhZ�i-�B��Џ���+ֲ�1����%���Mg�W!I�����-��7��s]�xʷMg�PS�X��B⫘@���PY-R��>i��t��r�1!�lq�"֊�oPh(��,)\�?^5A�,�n1a[�=�903^V��xд����`����L��لsV'�#�+KZ6L��1+�*4a��W��~+��.))B)�[�"Θb,����<��7��N�gLҺG곥X}LZI��D[���A��h��+|���3���k��x�s��߫��Hj��W_&q�xY�OB5P�����B���Jݷz�X�O����'�v���0����g����q9�$��E��Y1��4US�����|-��H�1��B-��b�T�}�r)��_����s6qV��j��Mj
KZ��c\��K�S�G��Ɔb�кAFR3a(�m���!�V��:�O<O�0&.?���b@�K^���!�.f�ZO=����������m#)�H���(��i(Wx�>Y�	� �EM	4g6�H���1���B��׺-/ka()U���J�=^���D��?�H9�@qJ���4�e
=�F
�j��)�� B}P�-b:���(&�x�����t1��z��#CM�!�����Y���REZ|���(�����&�Rn�m)�C��Aj��hV�i�MF�i��xߏBFO9}��p�PQL}sx���v��m��m�[۶հ14��&il۶��}����{]���~Μ93��g�$;ǲO�Ƕ<�'BP��m��<����(��ѱ0X7��\���6�u�(��!��Zg�.`�a����	�#��e;4F�'�-�r}̞��%���pT,��/4j��x�(o�����$����M��.�i��Hz����]wU��+��$!t{l�<��ۓ$r��d*˖q�d��� �������(�����p����pTH�����J�|�d֊f��I⮞�o�5��J�fK|r�C�ȳ��}�b�VfSt������&��#����$���Q�/����n
 H�+S�39R��0NA|�?C�\��0iq��g��.����h�͡h��ڂ�������4��;`��.!ҋ�ßB�D &�,�w�~��F��ߺ�����kL�D�!��:ȠL��H�w�Y-)[�´U�2���S��mzM^2��p���n��)�t
�|��4P���`�H�3y�28����q�0p<b��Di;�Jx�jH������O�+�AEf� �>UYE�WJ8zfd��*����S�o�g�yw��Y):�Y�_��YӼAu�$8�Xd1�T�H�M�sQ%pIGB�P@����A�u�������̽w��z��A1�Rù >�P�7 .P��K��:5k�lij��`�.a��A�=}pOa$��VO�U�����IU��o�}o���J�Js{�S�a�b����l�r.���;p���M��?">J`cE�y������Z!�BC���BK��2��_����kbש�|�.����`0�>���E&�oǘ@���Ɏ��O��'�g_J`��-sp���F�����\=�0���FE���/d���Άm�lZ�Pe�S]�e�W}:��Q�9d��}X5�qj���X>Cα�?�?M,���NW�L4 ��r���Bބ�s^fS��4����@��Y�V0�{$�O�*�OS?�J������c��V�&���U�`L߭J��bI���A��l`E�q�Tn�He).׆�*�D���TIm�����ҋUoA��E"��Z�Z�����n)�_�F�$��r1T=]آ,\�矬B2"�oD�)\�&��B-K;��S(#[�;��~���ms��D*W�T#��#��>j�ʨڎ�%P�����ZH�Ђ�P\�|���ѳr_簇������0L��pgS�)�EE0ʓN��^C�3e��.` ��-	��a�A�~R���z�?< {YB�O3�+9��X��')o��V@Q�H�a�Yb�;e���!�	�@��M�ϼ�o��O�R��=T��
��_|�D�8�|����	p'9��"��Z~Ʌ�q�͑Mz��_W2xc�}��R�\� Gs��� Ƈ�O�?�29U�i�0��.��1�Ig�����!Gŉ1U堜sF2Y)c�S����K�(�1����H�F����#�ɒ�P��� %_�'��tAMT�ՍP:]�Z#�Ĵ�;'��2��Y�o��P�5�2u�c�H.��R����z)r��蟡_�(�k�\+�ʡ�,��ґK�G��������r���,�*�rZ��|۴5ݵV,�o�]�𯉘؂��S&�aٮ2�&{Ootp��V��e����QwY����z�O���C�k�`�~��������	w�A��wC�G�?��V���	G�X��m%�k�a&�+˓��y�q��x��v�ߋ����%*��w��:.O
��s�ma���h�'tLQh?rҿGN��ߊ�����\�l�Ė�����U����F?<ʎ<��=�=�m��,�3p���lN�$��+�YE���E�%�>�;iX)w�D4�� u$	ޝ�{�:����'�4�r���eޅ�ک�S���g�h}?%'y��侽��d!�a��W��W�?�mK�8�l�+���{��
������`�h�_<�5,,(�]�0��GR�D<�*�I�����	%���J�*
!	~g��}��v�����7R�?��f,��}XT�?2��!��tg/�I6���j3/fv�7į���~>���\?�^l�m�~����$�	�5��1��Uh���G@�C����=r�aЋ鎚���kx���܆9�5	����+Bh}؞���\���\I��o��#+4��_��+��v0Д�lBn(�6Ig���G��"*���j~��,�.������0bO�Ӈ�(�:`�PD�T" W;(�{��
q�R�ZI���n2�4F����>��/��<�RL���QYm�NM���$Ѡ��G��N:��=?1���A|.j�S L͕a�;Ϡp"�˿����4��%V�&W������h������4��}�}o��^�	��It�_��<�"]��x�� �#?���ɖ��'1M��NIuD!?Skjf�($��aâ?��5�M3�zΔ�_Z�BF�O�hu q
X~?�|W��xp��`��K�;>�;m���9�-ٴ��o�c�+�?�TA�{Ca�oQ�-���N 	�W�ۓ%X���.�~q4�\Zt2^��*��P��kSX�)cu���-�?]�Q��lݲ�/�q��y�T�8�^�u�����6PL����@��f	��o(�|(7&�'��jԷ�(?�n�b���t^pi�֞�QM�V�}���aF[z�R�C0孴�=7_'�/`��h�G��5)�S�ӕ�9���jEnq$!8����.�v\��E�'�d�\_֘H+����BC3
K��묈��)�l�߸�h�C�C��]���<˲i �|ˋn̋XL��M����W��)'���]�N{Ã�A����?��G�FH��
�a��6���J%��3��>�~P.���U��gp�y��zB��9��'5�Hy��ݚ�S%���O$�����B���e,;�����%zDQ[6�^ �Z�'1�W�-��Xioׄ*�Ʊ�'丠f�IaCqpzb���ќ�*�O��	�b�*~�&��,�s���AmE�XN��rn\ǌ��t�i�_�����b�^Z��RM|t;���3>5Wj��A�e#�x&X�q��&�Dq�X�,Q͝�rM:f./u���'�)�U�%�hqP�V�cm��FTaC�ރ#�=�.�;dM�&���YԆ<5ѻ � n@��l����h�]޹ϸ��-.m�凵-�Ҕ�,_��}��r��a��{�"���]9�븕�Ce��5f�!#�7�_��QT�I?O+k伍�Lj����'�h*�Q�i�zY"��<��~�ke���4�BbR�B�
\��?jw��
#  pC�Q$#�������*Nu�H��'����9��(2��J��nq�2�=wwD�r�ƛ��*�<K��.�~���As��v{l�P�=�f���h���ɋڙ#��K�q�+��bo��2(y֎�U�A���'��|�u���+���gίz�%�g��f�x����+,P���h����a]�nD�͍�f�1��nŰ����G����a���VI��0�='+�E�'�)q>Ǯ�{F�%�ʚ����-%���zH�t �*�e����7Ɋ��
����#gO��C��h�,�I�y����z�bڗ;�3�a��6��s�l��	��qV� �צ�w'�����5JW*χ�3�P	��=�c�ٌ/	��#��=�?�Ŀ�XC��~j�=����Eō��0��yU����fgf���*�K�*�<��X3�]K�D��;�p�ƽl�Z��w��153*ş�k��S�!ྸ����СO�qlf.N�&.�F�F�Zlz*�SH�!G[�T. �SgJ+ר"��Z������I�!���$�v1
�䒤Y��=&#��U��,++����O��h=��f:�oigU7#��L+T�e����2S$�a��b���<����L��J��5�)��Ws��T�&B�s_���v��0�<��i�gRx���·��1n��i�M���08�̅)Ys���$8"��)��W����M�	�<��)l�fq�����S։�jMw]n���bJ�-��W�K����P,����O�?b�:�5���&�c��0�f�m[[H��*,��֧%XWt�a�[��'� G�*X-;�Ӿ\V�����d��.&J/	�����D�b����b�$c��V���:4��.�.f���K��[������*��q_�)DM�1�m�C��ωL�,����8A�P�n��$K��/���|������"+SeGx����P9�*U,�x~d.�B�t�\�<-A����6�3�+Ífs�L��Q~�q�~l_x@��h��0U��� �u5d}�/�&ņ��kL0��1aȂāC���#(��0s)�ݗSbpl��;::�9�F�D9&�}����R�.��蝗�1���C�r*�#���q��ӟ6�σ�M�/�rl���6C����o�-F`\�Q��Q�{�fzϒ��r,y0�N �&���������?���,ka��E��;�\�m�tf�tz�G��ji3}꯵c���"�����bI�;�3��M��K�(�2�s3�C3�H���lG�i���DLX�����r�8k\�o�e@{oe�$2��JGRy	�?{�/R��n���s3"7���j��`��A�^������6�At��i���s�N�u�f6��}��M|r�b��d���Wd#S��b��o������*l>:���DS�F��5$�nx'_<�v*�T뫧C�������J�*gA����$�9�Y��u�p]���R��خ�r�\��x���A���=(�&M���-�In6��P����� ��7�1�����v��o;<�h�����olǛ��%l2M�=t��K�Ru����L��z�i0�rY����x���u¤�(q��X�E]]���i�Q��;E�9��%dI�9���7n^l�%��0x�@3 kj�m_æ��j@���6�trx�˭���G�ω�Ǒ�,N0�p� �t�/�t2��o�T�+��fgW�qf�NI��q�Gp��:6��yLV�RǦ|��pdܼ��&`ս\-
t��<ǜ���N�w��)e8�eϦ~����SS���;/����
c�cb�u�W@�t���{����M}xB������uG���o�\��g]�CA�<\�(�⊈iqU��]fPx4�O�z(���.3�Q�ڼ����:�H�:׃����HB(�J%����Y���]�'���}��`C�d*@!�{rq�݇L��=��\�פ�Y��h��z�!Y�\���Tx��+��ĭR��{iYQ��nê�Sa8A�`�_���ZJe%-�C�ߧ�9bS̺UGT��;�����齇��ٚ���x/� �'rkD�>�1�"u#�q`9t.�w$��l*q�(uV*�
���� F��O1�ܧ����r/.�2���T[=�{�N�ܰC#;�\w���K���	 P (Q~)&;N|����ͱ���˅�4�JR�^㋍��4[>V�q��V҆�⼬�Ms߼������=+̆�������.K �m��p�B��y��SQ��#D|0̀	ŉk��:9;k�y�����z�����������~깰���y"��γr�~*Q4�Y]���jk�uT<�6�e��&�9��u1A�]H��j��-���P�I�9�5�͕��)0�a)�§�~�\���w��0���jqE����O��A�Z_:�ͼ�����Պ&�<8A (" %���ۜ���z�H�QT̪Q��C)#>�O���O�|ز�ls��A4�%��jK�r�Q^^��`���ǫ�����c�=�̂��ԙ�u����.������P��㲪��F���D��éFx�F-k��N�Qy�5�QB�W��hV���Qg�z�Ucc��l*C��EG��]��T������D���5��Y�������>'��<�V0�݃�1���X��ł��Y�a��&�25�[�[��1��M�@��1!��u�h��قP##<ѓ�G�'�p5��X������.y�	���,��֌�y��8:�=�A��� ����9�b�G9h��Y��S�����2ӧ7q=�ru��}E���/gM�[>K�m�Q��!|��,����~4���N�	�'80����m�k<�^����-�+��_!����nZ<�{��q�X���˷�}��-���#+�c��:��z��*�o�t����]��n�,��y�����Q�8��:���MFTl���ٶ���߮�^�3��|�Ӈ�YF���"��t���l�w��)�x�ۥځy������':v;�+�1��*9�_��5*����P[�U�LK�OM�1ZSx�e0b���4�Ni,���Fzz��W,��(�&���Z;��9�$�-��|R�a`|o�B�z�RZ����P�����]GbϜ>��Ի�:5�"��\������-]T��Y�|J�1�Y�q���<.-;,)�ͷ�����R_Ƕ�ځr����t������f�:���ʲi���ei ��~��s�RRٶl���|s�/�(�B7|�s�w^�ɡyb�O#�⏧	��	�{V���T��8���󶕋*�1+�o�'R�� �$��ۼ�Q(�b�L{����C|�]H����U����#?K��%S,ϕ�u�������Ϭ!�;�M�M�ڣ<��жx
 �`�����5�v�|άG�j�>����Q�7�m�C{X�����{Ql�����M4�*��U����xM��b;->����_i��ĖR7��/���_��m�Y�b�-�	z��Um;�o*�	+2���3<8�[C������g���N٤��i/��-� O�w�rW?m��O����:��K7E�K�3�=���%4� �Wy��E鿒��4O�8|�W��Fs}n�z���躝�=��I����D���DA���O�u�r�M�'�5�^��Pf��i��Ǻ��h����z�׆�?] �e�6<��#y�o[t��۹A0>�̩7��cѓ�x#�4����q��Z��W̯�����[�B�;+�}���V'd��O~�P���96Kmo��vzF�1"��o��Cp�AXQx �׉9��ᥓN_d������&f�%�~�@ɇ�^#�u��W|�?��%��s�����r��w(JT;��zpxT���0Џ���&�jH{/�؃�l���B��"Ύ��o����.��MCD"�]��U��U~o'�h�W^r�}�i��F�>���^
y�c�eU9�Ǳh�bVV�/h�/}�8/E�S[m-���q)�v|��Jp���J��*e�c�+S��t�Z���nq����%��|��`��y�L%<ڦˍ�5��%Q2��
���$���n欇�	!��a���ՠ�}V��6Ѻ��BAa�c���d�$V��3����5��ҭ#���R��z��" 4����aX.�V=v���&1�÷X<Yb�~bd����v�'��oN�o�k��WkHK??��=4���}iߑ'$Ҍ��Q}Ƥ�4��gs���p���4���e� � �`�.K:x/3��W��>�{+�c���e�=���a����峱��گ �kvh(S����'O�C1ڻ�bp'�
����$�o?���Ew �a�P+�;�g��N$�ňF��x�3�z���!�bV�{w����zCŚ��'��� ��Ey�	�����C���_2�4/�:�%�|����@c��t9e���["���%J��\�>��4���7���݂B�U�ޕ9ͻ|�=�C�ˋ����ي���r�?Ś��"Tj��f���g\ЉOT�8O�E��7m���[U�}>8 z�(I����[���������2"l�5@�ݰB�:����~�n�k+2��Q����#�e��c�}�Z�ʄ�ô����t=tI��6�'Fǁ��2
�bY�I����:��|H;��n��Tl��>zl��kxwY�ك=F�£ƥ���2��o��I���G$h� ��	�uK���s@\��|^a<
��O�nw�9�����_�)�����V�7v������2�ұ�Q���t a�\�
�ކ�Ā&t�E�G�?�GE"���Ϝ^}���E5���3����MA\��C8��R`��Ԕ�ˉ�W��^C��\��j��,B�`�d���3�ۤHD9>��^�=�q�f/mn�����/�$�P�o����_c}t����9�x�5���k�"�E�(�϶�'�g�u����	�n��o>�/��	��x�+�_w�5��
��C��f>W���*A*����c0�f1���sg�&�y��Ӈ/J�<ux�7���o�Q�a����G�5N��*x�B	ޢ��$"�J�O[x��)s�@�����&a7���b�}��5�;;��1��ǭ�i
�M�n�Fߖ��g���4K����znp��`��2�7@�o���]�!��"r�ہ���s��n5����f%�	8L �C3��+�To��_I�[޻����!��R����rR�Y���Q6I:�Jr���)<���
FG�JKbx��0c��鐜�̑���m"'�ǤF�w�]|l����s�?���	��Dρ�G�1�l�_޹�#D?ym���t���2	|�V/|�üNo��<F�>��^�Q�7�BPN�3O�i����3/uUM�r��K�'��D�$�*.����H���/�/��_j�g��K ڏ�&d0 ��I��G��8�P�g!��nJ�������w&1 �՞w���M��]}R� ��gM`�[7����A������6�p=B��Xc4b����uܱ�y=߼��fC<ktb9�Px7(���̱Q`T
UGy;k��C=��}��B�Ná����hVYȊ?��3�������G{����4��M�M�h�Dw��Yp�f���v�lwlu��B���引����<�W$L�W"A���1��=�.L�G��D�����`jB;��#��AH���>�X:�E\H��X��a�!P �'�׫��t��gX��	�M���0�@> ��e�N���F�����N�\�h�$��U>s������r��7��
��g����/��y����Vg����j�M�Go����߯����v��i�d�<_����Bq���q����J��!6��|�$��b�&���{������}~���W�Y�:����������m�a�Jn��G��}n�������[%ֵ����r��A�nC
���Cf���>�#��������-��2���>ܲ��dF��D=}�(t����o�U;�_[��C��-(��+^>-��ͷW΢�왺QokՇ��Z��p�I���+�ٕ��2e�EH^�������Q�
�
�?�C��m��P�� h��\A�HHA��̖�f��~�Ա���Įf:Fx4І��k1\DO��q�*��ȥ�E��h ���)4�{k
���x@�6db2���i�\O-����L'���P��';��������D{5."��;[�y*�����2�� ��W��4���'��e��}j_ε��n�-��C�|��q�h��k�B�we;9��o��c���?�����\@����$P�	�K7�wt�q8J�V�{�b1^��!��m����It.�)K���=�)�iը�"��?��_ae�	L�y:������ �K;�fBpC wo��q��W�T��W�- �6tx�	����v}l|��)u��Z!nZ�o#awxgŋ�l�J|'G��fd抻z7��&ք}ٽ��σ8���Y���@��j&>V*�Cx :�n�>�I.8䐅��2���g�z|݌wg�v�m�?F�=I�\��D�{�d1�� Dg �Į�$����yۛ~*����V�W��$�]BL�-`k���وy�/�l�Y���������w4�'��/�s"�ڷ��v����ᗟIf<�q
D��,�a5��9a�ȴYQO���.}f�pZY{jJ�o�s=����#����禌V��|�1
s<���K_�����~0�ʿ#�}�P��S�(:� ��Ar�����i�'�
{�R�HCQm>�&N�Gͤ�mL����O}�4.̓� ?	���B�P5x�uZ0�7	��`f"�ӆtO�c�s��u������id3O�=q�͟�=��} ���	���j`
�9Ir~1�^�4�=tN��Hv�����@��0�m���s�u>�þ���]|^���j��6욹g�o!�	�i?�<��վc���^�n�8�%��A_:\;y��M9�pqb�%"L3P���y�����U1��^�:�idEH7H(�8m������L0y�����%4zR�MȞ��\�R
�j����u����f�N��g�0�]j�'�k����N[''��T����53�˪q�5��S)1��uE�Oo*f�m\<e�c�}Τt��,s\`9�cGJ^�"���~�1��C�ZoK �#�K�g���;��8���No݁
#�b�G���qq;��E�D���7AT�F�SN��dV�h�>ސC
2􏃕�U�m���^�����}.q��b8��s�a���[�$���ؙ5L��p�B ��~t���O� �0�ND�
���h���L�7P{�p�z�y���=`�Xb�[��L�-.X�P՜!������� σcAH���C)�(���O+���
Ry'��� 1��H�+;7 �p��:�A���%8����ɰeW�b29����/��!_cvW$3���7}���h1��N1vnb����/A��^CoF���p��٨�x�@/3��=֐;ӠC?	iP�pnU�!nr�H������}vU���S\$0b�������`�z������	ɶ�RH���-������SzImU��3����������^��J�"S@FN@���m� |���j�3��r��H�mX.�Y��}�j��+z��Srx�v�\���Q���X� ���@�x��Kb�7��$���Ԋ��6SU!ڃP�����q�Չem\WF�!iN�Y��%;�L��*%��qu6^�8~24��ӳy��T�F��i�ҋȄ�\S�YN�]���Dj7i�*�il>`=ņG�3�u`K	=�/���p�ol�A�+�q��>���ScLF��'�K���*�����>��"��l�sp��e���^���5Ga�o�!JF�J�)�7�gP����|����`-�ڔ�{+
�?����Ç�A�����R�ǀ"�q��
��{_ ���=�&<���{���M�I�&��F˟�]��FTl\�;���$}8�p�5~���(�tt����:�)pq�1���[��1	���wQ'�_��c����m]��u57��u7��NZar��\��d�"��J���3�͋���0��ͻ��{G�sm�!s"D[��"���/B�(8$&�嵣���y˹�\�k]�q�<I�Pxz̨����y�=�| ��u�`�����G��4w�R,+*6���׉�q5E��������d��V'(�L�(@Y��������{���C�����a�1��;����!���?C�Y���eCn�~i��4�> �BF�*ۉ��I��z�Y�T�Jw/u�&gR|9a��x��Dâ�bٺ��dX��#��� �K:��L�U�����]t�9��\��כ��)��o�D��]��V��}TX]W�H��LZ5�pf�Clb�}��W{��"�V7.���h{�@E�xMނ�|pQ�۵���)�at_��L+�lZ����і!�3�l��G�;P���´�)��9u��{휧����'�l�#�O����Z��覀�β���u�q���뚑�T�Eǉ���Q��!�ެ������t��qދv*]��\F���^��x��6Э4�-� �gdL��h/(�����XG�F��w<xk�TK�T�-���:,�l���ڞ�F�P�����5�?9�a"4Y�8^(��v&%v��~��:��8�������MY�(���h��,7�4��	*t��l�"Ҫ9v6���,�&#[�N�7�2,�-����em2��AWF�8�,�a�q��b:,.�'�sU`^͞>L�g��銟�̆(,�t[���+���y>�&��}��1�rc�aρ$f��1� �4#�s��@�id���3S��C��$C�����`8��r�%V�Cޝ�p�[J�����? �0u�׵�'pC���8���^I �<"G�K��
]t�G2��qp�ų[�V`J,�ݼ�>W�ȓ�,�H��$JN&���q��i��o�ՁjO���	�z�-מ����YEX��/�+�}�e�CC��b�Թ!���\�>��x��9����9��vF�	�F�iK��C��&���o��9ہH�rT�}1��½��;d�#�s3a��FsHW�^�7����D9%����d���jSH�ĸ�cc�6�M?$P�����:d�\�`w�N�"JQ��8 �� UVvא?Gr���ǣ�<Yy~	���?�P��mz�)�;�ғ���L^�a[���D��Z�E�F;g���HI#��u"uX3-���#�{r�yt;s���J��Ī�@�m'{sSz��%���p����l�Zw߼�Z���aAu�:�O\����?��E� ]F���:��c��-�)�{ �q��zEV���7+O�y�"��1�@����ke?�-ċ���Rv��q�GH�ĒQ�w��Fcm
 ���_�ϯȕJ�1nX(ٽ�幖��h��`X�uz���#��D����S
i������D'�Q��G�"ߔ0��"�to���{4#��l��_���2�-�C��|hyy�xTƸ����3.�8ʻU��^:~x[�j�0� r�ͩ�S��y�O�.�mPҴRO�!9E������o��{`��O��Oy!9�x~0��[>�U��o|���K���+��ZBs^N^�H��9��F%��!$˒�&/2�g?~�/?��#k��޳���f�J���No���0%�6Sy�8��vkF.Q%?�̥~9̩�/�zh���`��YA�-E�����&�B�C��
n�0X�o"b�(��7���ʗd�<P�PRq�� 0�W����Z��ӊ>�^v�x��bߠ�Re�~�Jn43���m����Pb1��C�=PxN�AHx��Pe
	
9T�����Z��Y�U� �`�dD7:��Kk�8�(E�`R��s	��ĠJ;�D�%lL極��>���5�;UĊ]��_L�$W`(*��z#4�,����\��!SN����K��r��C[ѧ�f�0㗌����#"=z}�Y��yºU_�(2s��6��"�/T�c�4ULs/���j<�E�1B^m���^c�c'x8�
����u��ͣq̌˗Z,����xao���>�'S��ފ3���s�,��V6�@��xC���e�F��z�'����1F������&��x�
�^�z�h��	�4��� �/ʝ[o�dO�ZA#{�̨KI2��$$H�}�%Vu�1�0��_KC��LR��[� �xo��� cppN2v�|�������-fh"o&�;��X�m���jJ:>L=�/����l��d����n��x���UE��	[0	7���Ҹ�<?3����BP�=��+`f��,������)�M'l%_���d�>\Q���n1�;���&�*֩`����Rگ"��R���d�g�S�B��W���^uòU@�
�ax��<��d2v�p��Z��$Уo>:��)	O�7�Dwi�Nk�c~���t�
��^&����)q�B��I��2v�
�OI�(z�m���B��on���X��8c�֠[f�4d(f�<�n�DE�n�!3�hΜ��.?=��������y.O����Vz�X㕙
�On\Q�S8kc<�}/nB�D �����K�W?�/B�uO�#0���֊�(?cG���g����\�^{������<�����=�S���~\"p$���p�ݞD��
�|fL�	 �����?{�a.�r��.z��?��cu��x��l�n*��Cb���Bp����@QE�� "��""0��_��7H��0E�P*"O�����6��n��7cNf�SS@3��9�O�{]���ۂ�����G����!�s
�}y;�D� ����`�iU:-,�y��,W;��n���X&q�3z_�����{A��w��lV�����bA��U�v�3z��'�r�6�W� A6T��M��s@�"°XF$��w�ɓP� ���������yz�W���eO�7���l�3�/�f3J�>Mm *���� ��J���:u�􊰗�֞݉���g��eX�s�}���3�gqI����xy}�l�r]�;�eSĲQ�Z�O�ϵ9~��í��{Yca��ī�s�~6��ѕ,����v
�ȃv{9s�p�I�M{���&��BU��@,(�'q����v���mu(\f�>2%-���=��>�����^'�%���Wh�(��;���X����b�k�y���a�B'��וC��N��HH�6���]����vt�Eg,iF-������^kh���9�x����/�Ըlt�0�:E�B~:��:Y���]X��}�@6z��zڑ����ˆ:Y��^Az�b{Kx�gĻ:�[�Mϳ��!Kr�ZL��D'|�^�#��&�w�A>/�?��tD��yܡ�������?)J�db"q$�\;w�`�^h�w: ��<TH
�s�Ԅ���\�P�R=9���;'�}����̩��q���~����r��L)��L;f�7b��ջZ��@�`�ФŅ���:_�G�&I�n����ґ�h|�^'��po����'^2L��0Z[��gnw�VD�9���c;���/��јVJ���;8=sNy@���/\��qRP�#��i�XV�:6mo��`�fy�w�?�&b����J�.n�k���� �p/���C�޹l!J+uc�8�sW<��A��3�a��#�S�BWLE��P�R���������g�^l#�~����fj��כYK(&�8�-��@�⾛K���#�ծy9�a�-��'��ש7k�&о�Ćg2�\��_g��J���6�|6[<�7��$�j�����\�(`�`��73Gkg̲Œbѻ�j�q_,�z2��}�v��ڻ�"r�Đ���P~!@����x Թ_�J[�֧���XGרo��B9��8�I�0��(�Y t6�IP=_�M�Y��@z%�f���JA�\�Ԩ��\�6a�-;��j������:$�I6�]=O�Oxƺ���`M��F��RA����bv˴�5�spFp��ǻ����<g�Ύ��7�*��(�맦X�?جe�t���խK.ðCð���U��T,�Q�3�r����wP:l���ٴW��8���)]��	S��Ճ�:� �AHV�'(ͮTvA��2ܽ��%�����0=~88]R�nG���H6�8�Q><�
~��A|>;_���&Lt�ؓ��;KS�ؼ�y�N��O���S���"�W���[;r�P淣�ƿA�ζ��^�
�"��b�a��S���'?����'��A��{;��U' "�o�4K�e�)�B"���������˥QL�=.b�J���m���U\&{��-c~�����F+U}�;^�!�ҟ�=��qej�%���w��S�`	��U	6�@�ƾ)֩�n�$��i<4W2�uC;dv\�E�_��3 ��<�H&�}�<���M_jS�u�!�����>������.�4�L�.�9�����
�(���v#a���L_�i\pd��o�O��j�C�(�H�Pfð�X:�}Mm^d�w�<N�|�zi�FPW�m������@�L�;5�
�Y�������}�~Y��wJn�����F5�Ĕ���Șih~2pw�n�'K����|��w�Q���ꐽP����tń��q�S��ЌDP�����B_��#��жR�J*dx�NF�	N��c���!Z�m��N� �Jny���8��L�N{��7	h��J�P�6�q 	�]	���r@گU��0I�{���{<���/	Y"W�p��kw�s\�B�k�C�7�bI���c�'N	w�H��RB�l�=^�U�^5�ajQE��G�M�Z����gg��I��
��*۔�#�����L�2�?l#ŉ�0������C#��:ա����JX�W��g;�H��@^�|�U�3d%㨷��U����A����=�����Q(�dc&ܫW���}�p����c]�m�H�� ����O^N T�ut@��$H$����a��x�ك�\�9f����{vJa�]y�>+���Pr�D:�AaZP��߼̗�!���>���@�֐���t�ny�``O�4]eX]�����Nqww�).��-�]��[J�-�(��w�\ny���N�̞-묽�3k<��)�kl춧Xf�2
޹�j2������_F�ޫ|@�	ÖQ�
c�nt��G�]��3����Q�I�,��>�!��m�G!(0�������Q�5XN�Z�w����x蓲�I1s6Ό�3��H�B��?&��k.��O(��RZ�F`���_��0�b9���E���Xf����~�)�����V�2�ݒ�-�'㸯1���a��!���͓�T���p�����F"��^��N�����&\��Am�O.:�`�<�J
q�[m�թ-W�$;��"*H.��{�O�mH���@Ҭ/~^o�:k!�l��M!��jG����a]6��7>��i!w�&ҹ����W'�QR���	M� �p���k�.OLŝ�a+W�¥�Y�z�¾�e�m�Z1[L*�N����s'~<A�ki�gJ�O��#����Q��XIr��m�rrٔ���*�G��GD��z�*����y�U�Ê�w��}���"N-�t��o+�V+o���ա�c+N#3i���䔕�bi��T���o&H�S�~�N��w��!1���l���Ŕ^���6x�g���;E��������ڻI���oe<\����1�x�M��J�HH��]=ր��>%�a�p�������a��6�9�����);;�A���e����Vun��g�kĝ���,B��I�}�M��j�O��D�X;q��g(�� �U+,$i�������pe��hq���_��X��?[N��yxD����h���������(y��gj� f����0O�&���t��7|���|=�9.�Y6��ٴ���2�u@�`~K��K8��JN
�i�c��uU�٪�g�Q���|��R�������������x�1�-$����F�>�g�Ӗ`�B��"�"� I����[�F�9h��G�V�Ճ���E�l���f�J:y�P�u�l�<9p�v���يr�JƷ❇�^�wx�[���}b ��}������>�90��8=#Y���ć����h���` S|ОR.�d�G?�^�Nr9mx�15s������/��q�U�sv��ԥ���E'�1��#��2���[Z���Η�Y�y���&U$�$U�)�O/�3nk޿���R�@2� gK�_��ww��M--���ַ�:l��炎��(�yZ̩�����ګ0�ύOăSa�w��ܮRW\��-G 9�$�Vj�|�uQM����b�����A?��(��6b�+�n����oj�Z�G:�'Һ�JG~�"Q�%��=��Ձ�r���.��|�S�'։֭���o�����u���B�&V�vw�SJNN�ǓwG�?p`�c���[��ޜwN����t�ca����I�ַآ�5{֣F�]�	����'���8�|/JF��?�O�%H"���0���i �ؿOs��M�;��=�ìa�Jף,kMɘ�z	h��˩�������ĶW���=}{
��<�%���EHp	����I#[Z͋�~����7ɨ�zn&_��������t��ć
��f���O(|� )f1��b��ˎ��Gm#���Ll&K���`�dXpQKc'=ޚ|�f&ݹߨ����#� ��ݭ�zx���;g�>�@��1A���[�5�=�*���g�4l�A�w��{��z � ?W�} �2C�T=k��b�r�>MB�S���ܥ����/��E����z���t�}	�8���G�2G�s �=3�����{H#r�nn��%c��Y0.L]v/�o֠F��@/�a��������;YD��V� �ܖ.9�p�y��E����3#�����G���ʼ����̛��nb%�E۩����3("MX�5\�Q\��%7D��b2�S��R0�` v��5S��O�R�M�x�
�Cz:��{����P���.岙�B�[�k��~N_^�^�%W�\>+�Hַ�g�g��
�6ZEm:��蛡�V�<x�xm���Ns��I�w�hӊ6�ٮXvLǄܮ�_7��Ю�F0�~��+�}��n��7�r�>�,C�_���4��xq���#T�����V(��דL-��اm঳�∱���ӋAI�=6@*p�i�e��������.�c��Y�z)�lG�+������;c��$�����Q�o]��(2��$q?��������L0�,�d��Jr�n�,����8��9ԺH�B��JNj���]uU��9TZcq��8Y��P������`W½UZeO��W1z���O����݀B�Ap����`01)�j��6�iQސ�Kq,�2HN��vӕ�$�i6�ʺ�;p�b�Bk�j50�v��K��VX8�Iy�IЋ�JLy���({$
,}f~�+|'�v�%1�>���m�f��6$jLH0d fk�'�Вx<=��N$Y��Q�����s�n��L��ʐ��C��xH�L)����|�͊n���U�R�nM'6�9�Pb8~�	��w-�8m��6y��ʼ��J=����bi��s�C��D�H��c���TK�K�J��˃|K��N���c���C7��i��^���f?p��:0���q�.�� ����`�'�aɸ�x�e�ɪF�]�h[
��
o�a���'�k���n�Ѧa����2(��Mm&<��ƓI����fC�=�����(<�A�����]	T_���5�~���(����+�C����K�롍m�ۼ�d�3G!8J�P'�T��B�8��>@A7��$��XM>��7Yǂ��W^Q���&��c�Ky�d ��������Oڷ��cdo��;��}�ۂ��P��5b+A,�%c�,$*է��|�m�@�3��#yO¿l-�wY%��H�����M�drj�rҐOɲTs�mz��Ý�ѐP�wUw�M����J�g��]���ʾA�O�ߟ�	�)B��5����m�Y�Lsi1�,��O�qr?%2U+T4y�_/�M�w~a�`SO\zTYV�QH%D�k�dq��l>��*������ޱ��2(V�(�@w#^�|�u�����I��8�>\�d.��'}���(�Q��E�j��Ĵ��e��^��N&f���3�~.��s���G�}����e����[�3���]L�<�t7Fj}=�.JRF�h_��8��4��>���m[S�ͺduvN��z!��h0�օ�@#�S�oϱ-��ފƿ���Ӿ�rsS�9��]6����S��@:�! �~�����V|���N�d���@���ï��_WS�l�jh�;��joB�dld�.:<���n��Y�kP�:��!����d��q<Eٞ<P�{�8A;A�.��ӏ���	F��|E:Z��cC������C�n��Җ׺�Ҥ��~OV�,~\v����α�Q���b�ᠻW\p ��f�oF+[���.N-L%M�ݤT��;yN��F|1vǓӷҎ:��<�e]ә�S��~`�{[�Z� �o�����Z/��R��;��9��Ɋ9�/���(��\��kR�<��3p�.�����/dq���Hd3O0�PF=,�4�J�4��$�l�z�_&4*G�Ǉ�Bo�ۇ�3ya�ӥ[��??��3A���k��E�t?X�Q4�O�Խ]����pD`# ��j(��q������F���̵�ʉ�(g�o1U�x�MM��/��i��J��ױ�7&�l������.t�X�j�3R����<��a���JJ�j-�[Ucdv�8]�?25/�����,���������}e�b?G�_c��W��*f�;�>4��z�I�.~4T��v�q￪�b�e�O��9��I>+����h_g������F������Q�0����4�6hv���v������f�
���k��O0���`C��A&Q�u$�5�]$i�bW��?�LE-NײY��VeHK	�3��S�Uȓ�{�o�짒�T��ze�p����}mL=7�V���*ǰ�t��q\l��J�fy��� b�.\S��'~��?�E
oq^�栬�9��E�~��MN��,��3J������N�k�#�N�h�_Z<�������B�Z(NL�<W�S��ր`CuQ�ip�Z!�V�+��[D�Z�W�rQl%�!K��n*SE��t<^�F�a�w9�|��Ƕk�&���X�n�!|�~��Ǟ.J�����ˇ���
���{P�8���0��I����$�6K]cKM�q^��Y&�swAr�v��+���E��-�SS�X��v���������~t�c�̲��o�L��$���������2(�o8�!j�����PF��^��ę��P�p��&m�S�@����`�)�~	�D-�B7l�8<�Y�Ո��ҭܖ��?���p��R��I7*�'s�[o�mۮ���k1��U&`8^H%�Ob �\���r��N�S^̆9�$��v�;C�U��K�����~Z��d͏�'+O��x���,��������	�B�q�Ѵk�X��s�e�$�ɓ����ݖ���ߖ��Z��������aod���amfX�m��"��Fq��W*F���<��]����0�s���r�na����U�z�
O�v �y����+���Z�: �5���F�5Zn���(��m>eI�����9�p�<%ݣs	�m��y@LQ˅�� �.����R)W=�5�}	���/���onsj������ũ�$3o��²H��÷�~KE"d�!� �j��^rI ���9@�D6�(WulO,i�l=�i��\?W��8���w�4�G?��z�#�L��' ���?f/1؃Rᝋ�(HK�)�����U��̗�/���97@5^�}����;�^��!����LAuiU1�}\Mm����^5��QB(�%�+IQ��Z����iG����3)��K��T��de��_�|fC4h�5�?���Z��b���٫��V���[���� ��:��㥝{���z�jt4��Ml'cl�ʐ�Y�%&�R`��2�Y�g��؋�T���������m�R~��W-�p
Q�4z����EA�>@�~G.'�ڿ�::-�mGH�a1}���:�̞�����֮z��F�¾���[���{i��N}`�R0����A���:�v&7��M�O ������'���!�F��3��g��>�{]�@��q������J( �b�N�Y���O�����������[P4�@w�S\����;�Ary�0��Hv�����o��,�䃷O�o����5���A��rJ�n�'Nk����jn���+]8N���{�1W������NE'-���ݎ4��Ү�=pk{>�g���U6���	�P��XnNb�*8�G��{�����*A���L������<#tt=Ӓ�T�疰_�T�KJKƶvv���d��5��q5��W����j�=�3��:WvWe8�d�
;�Tҷ�]}wa����q/x�|�����#�w�fv0?��,�D78�M�3I�^����蝉g��v�+���_+.�r���+��m�-@j#���o,�T)�
�8�4�����@�E0�▐�6ͨ��C��w�Ԭ�;_m۽{���..�z�J��J�X��j35�\bs�P�ؑ�ԧ�ޕ��U��U���@�hJ3���"n}� �X�QB���۝e$�c�z�2[6��J<fv�,_lK�Q������9٥@揷���u�n��n���Xe���H���Vs�����c������m;�N<V���2EV���Ml��Ė�����+b��vJ�;�l��!4L>�����ɣm��Ʌ�;;�[-�:�������[���� �s����rJ����-��i���跳�����%�� S��=6�C�D���3Φ�ȕ�mJ�F�c�C����z���b�ǲ0�xNЙhR���K��D�+������b���nRn5��'w5s&2w�2��}��Z5�Y�Sz��:����%c9E|q���WŶ��%vi�������L�/$
kY�� r�d�|76V�8��\�:��H�rݰ*˕0c�:�n�
4��k�m��ψɯ�+�IP���}��s��M)8!��.���I�'��?�*����6�e�!���<L�M�R���d#�#����_����p��01#�:�����5n-�		JE�-�O��{�y5*���ϼ��\�(d��D�Pr�X�!M�3֯�л���B2��Az�9���o���13�L]]����A͗Jr�k�0�,=�H:'w][�ۼ��;����Im�e���� ��R|#X_Zpa�0�8��z���Nn �a�����wCy���0T��)�Z~�)+zO�zVɿ�E�œYyI����� z��v��t��[�k�@���9��C�(:�Pt!��o+�k'§���_5��\<T��Dχ����5�����Wr�P�!̽Q<L���(J&x�l2�m����
�����Bl?\�H��tn�@�0gTn�PG���<ex��g�ҥ��9XҦ?�K�B��k��a5R�T#�I��j��}��H0{���B~4'.�rG^�$��?�i�խ^(4���opt�<+��s�r�lh���	����r�ɡ4�p�뇻xCM�WV�u��hr�D%B�
��>��:������$Y_���Mǒ2YEBr���,����c���\
�[�C�t�a�>CE��i�P\c!�sW%�/���#�rTr,�W!����<�ij�G���ߘ���Ȯ�FY�'(9���b?�\]��=j��#��/Ó��������҄���G�kFN��!�7�WK��9��-,�5o���m�0<�>�c�v�*�%,�=��Pe)؍��Uy��g <����$�SsjS����g�\�̴R�tGs~3�c:�!}]qůȹ�q}J��u2���2��7z���,o�\/!�� 0�9�<þϸ�t:7�δ�&�o�����Lڏ}��VYޘ4�SܖHXk
a8k�4�-��HT	#���(	��e;w��S�=}�X��2~�?
��v�2߭����6������O�0O�2���?��-��|�C��P�J�e��d5%�x�O�>[ĮS������Ԅ�)�%""�j�-TءMΨ��C ���ظZ<�$�m��X��g��S���L��Iȏ#^L�[1�
@r��Z�����2�8��X�?�x1�<Q��.D蜺+(S?yh�C)����l��T��]�e-���b	t�m&��y���U��P$��s�������g�>g��k��MN&�����w�o֘��)���V
Wn��|Ֆ��1��G�1�q2rq�����^9���xϧ;׺؛&�{7�?ٞc��0���[}{/Z�I�H�	׼qU�i��p��Z:�H"�:�w�ѫ�(�D�y)�U��B��j�X�}����b)V���L�����d�xË�[A
��� ��ۡ%�{Ç4$von�i1�����F[L�����~"	��C6��iG�p�~]�&�}!�f�8��z�י)~b~excs!�ޕZa�0�=��(
[�e�Yj��@`�X�`d~إ�����hX�G2s�I�2���uFMph��G�벏hd�il}��&Ϫ�H<]q [B��ǉ3�ǽ��Lp�R�8���MJ��J������U�����tޡvY��kxw����,dcT�����=mS	Z�)����?�m�$ �������7������xO8�]g%tN�)Ո,h�.I�!M�dP!���xhK���C���i6���/�`i\�ݚ1\��ݠv�~�M��2�?���L+:-�ΙQ]J+� wCR��܄v>����"���˽Q�G�%�3�B���MN+^���u�n�A���d^��� z�P������ F�x��4/�$���[�K���:�|��F}�Y�do;��\�}� �߱�xm���,2�띁��;[Љק	���i[��f�Z�6�����z�&���X�*
Q��s׼��.4!�h87S	�l��/U~;tTY_Q�QaR2���3��x_K�Hw��`��1g�
���C�k�آ�D�iy[_y&��喐�U���H6�K���T�zY(V��l$�пv��tJ]���.
Ҙ��<��a��H�n�M?܀��$����c�t?�	w��C�	]5V�<}-0�������0FOgzp��m[����z`��Ʒ�wN�<&楻
�.0k�Lz��z�Ѽ�G|b�Tt��Aj0)��9y�A��#��|��e'k����:�������~��z4��@�g�@�b�����I+n^h�)�#�:.�bk��)���<�9�>��%��!W�Zpn��g����%���q�nb���[��^�ś��󰐓n4N���WM���b�3�*ecG�G�T$w<Y~W���UV�d��~�K)���ܴ�$��3��P��с�L�|6���D$��^���n�٢1q���P<bq�iF�9E�5�x1	�[��|hy�.c4�s:��*�����R$�����M�KhU�V�ݛ�UG�E%��Lk�	��'f�Uػ����3�9�ߣ��K?�Z��XOR��n1��@q��:�vV����kѫ̊�:��4���uE&���P�]����+�<�{��.���9/"�0�@��Ð����{�K����MoS���@��1n���H�c���m8m�%��.O��aá%�2������}��CE�)|��߿�?U�~�N~��,��?�r��8��k�m��XլPV���[���Nv�/���h_���_�c-L���s����^�Г"l�M�W�E�޳���j�"Rf!Af��j��!�_�2�5r ��ǉ�74����C�Y[�4��
��Z�/��D����Z����<�&�9d�`M/[�;�\7����%�f���1xv00��H�w]{�]l^�3��^W;�x����C��-�u��=W�X~R��[���X��Ô����sN�C��4����/uO�����_�P��o_�iߜ�HU��U��ӏ���[s	�m���:�K�%�@f�W[��H\�H.i�� ���������HohAk�Y��KK-�'�8��l3CR�/��ʳ����0�z Fq1��v�)@b�+2�G<s�aE%��I���zY�Vc)/�gS��s�c�����z�Yߘ;Щ�樂Cr��|��Y#q�>��M��}f7k�q��T�R=��,](�eyiL?O������^1/�n��T.b�f�'��C��w���S���鿰�����o�|��1W�jI��`6ń�)����;P]h�qb����zSiB�ju�ׄ�����,�?ޜ���	[�O���fT5�!�8O�5�����Q�h�	1�`�S+�0�wE=^S�^R��}����v� �	��C(��2$��!uM�ț��}��o�gI��m=p=_�6��m��x��H��7�>�Llb���\�T2UƉh!擉y"����s�ջ@)��=x��7��.�ď&P%EO�v��_'
Q����a��K<X��,T�("��>�d<�_'�ʤ4�����|�p���W9�;���y�����!��6@��S����IF���0�x�J�4f�׎ӄ��Ϧ񒹮:_�,*
�Cw�Y��K�r�4i���������Ź�l�[��kcǀ�a�.J';�U���yH��8T5o_l��e.h�s�p�>8Z`y_��*{�Nx������x�žmP@*�RAjD�G �IRx��M`~G�)p�Qz�Kxm�"
���b$^��+y]��� :����"nG�=�5vn�m����8�68�"��SB�&���i�w@+\H��-���Q�La�E��R�,gJԮ�;�R����)	�*ת��z�*��F�;'��ϽDc�}�]G�I���P��^�KAH����:J�!����}I*FM�}�*@�a��Y�{b�7��0� ��$��0O�٧-�N�wGxwr}�����4�fj|�A�Ms{�Y��=�.�`��΀<�[���i�I���,�~� ���7cj�m���?�f:�'*��$���p(I�Q�}�_\h�|vҎ�gP����A���A������>!~k�2�wTV����r��#'Ьǥ+"���qFr��-�?���./J�_��E�n���r���#v��iZ�)3�Z��It�th���B�4FB��ߴ4�K�7�N�Wp��.���i-�_+6���<��G�Uņ�^'z3�C�l��j9�ȓ,��
 �U�(���m�X@����oWWt/�~��OSM&�%H\���T��1���-/��8/�o�^�L�$����j�k��R��,Oqlre�Vg���X�s��ZG0^+��s.:B�~R�-�7M�LuN�s�����ֹF.��]�h��c�dt�0臒�)��
�0A��d0��6?�S�\s)��޸�m_���Ee�u>�Y���E�~�uK��c�4���=ql�Z�-dZ�|���\.�DG/�Jp��e�sE�}��6hr�-f�s�iu�9Gr��.I�o�4�9ȡ
4϶}�u�j���q�u��Q�6��w2�u��x�$�ն��H�h^�=.d�z�M��HB��6�^���N��.]�yF�If��M)�m'�&�B)*Y���(ݚ�)~K�=�/k*a�v����Q�����3@�'P>�&̦�j����,��7���Y�*
�?��ڐq�1V�-ȓ,�t���3�XY��:L'Z�aHcrS
l���&a�J[�@�g�{��r.]�Cy�L$z4<'(��ncܲ^x+
��K��I�|��[mԳ��/kZNjPy�Փ�J3� �/폀��o�[�;1�����Q*�	������U���oj^�H���Q�Wϰ�ݗf��+��=E/����=�2,4؇�Q��Y2ݰ�o\�d��X�c�2OA�OS���l��t��M��Q!-fۼ^컪�櫓qA�p�"�^0=��p��v�:Q���HJ ,�͔���Y*br��<RJ�פ?K�������Z+o�O�K�b"kc6Q4�\���͈Bo���J�=uQ=I3�So}����m_��&QC �_}�	#�^��g|�tiW@m��6w�
"��-��*/�P~��m��-Ս��o�#�ƾ%�z����An�����V=��]���!�M�O�j=zK��8��Ar*��M��/�Z��])-	K�2(fk��۠�"�u�$-Ӫ�:�d|vq���w�gr�|��ᚣ?�h�:��!/9��y�m�f#�J^���\
�F��&���֐c��g�J��*���u�Tϋ�ſ��)�?��*=�O�S���L���F<S��3}'��I�������Kk���������NZ�	�0����W	��6��m��S"Z��ζ�/��W�BWGT�`�x�g�C���כQ������T���k���Z�w�^Z���y�}/5߿�>��*.V�o�)�+͙2�QA�S:>N�+��G��%j�sp�����P�a8Q�7�lo�ZEP��������Ѩ� ��̿;����l=a{�*�'�R ��.�/�3��%]�`"�f�9�V����s���s�z�nL{Т��y'�t��P���>������W�����J����X�0L�]X-�����8[�C%'ϧ?4�D��O��r�nd�a��a�Wss��N�O�ڞ��3c��(�dq(Q�����Xئ�҅�|x7B�ǰQ�����T�ڪ�?�ؖ�������\g�����hvDhD��C�
�⼨��
���z��{��	��K�ی�gU�!ɇ����9��:S_	��&h�zԊ_��ϗ�R�MV����F,��$��f��ς�+&�#�������r3�1V?��'�'��Nӝx�$�|b���+������}��+=�,T2t1�v%�i
z�IG*e�����*�3���g���i��&��H��W�M�N�ƨ����_/�:d
ߏ�	�1G�8�n��1�Dd��j�(�n����w1�u�3�z4��AM�A����6h�����~�v0�t��8�(��ħ�hk�^Ϗ]?�%���_ϐit.'}5{h8�+Oa�£>��Q���ФN�Uu3����κw�~����Ӗ�
꾴� �l,�"Y�<��))�i�rq b[s3����_�OA��g�����i�%1^M'�A'睘�jWNw�!���:L���7P����琶��V��߿w��5��<���v����B�ʬGٮl9�\1��_��x����,cZ���q2��8׎�����}�J�{9I��U\�]�|{k��64��Ҟ�ߠSL�\Β~yi͈��0f��/��)��v]x�"�I�59ev�~������S�P�w��ʈ�����H�Ӓk��i��#4����nQ^��&b������"�2�0��Ʀf���o�� na�(��������G�Y��mv$<�|�__�v�oN7Uy��X��	����Dn�|KWg~���0?�;�*7b�2�i�$�������$���<՚� ���P����v�`hc��	 �O�jn��~��{ef��(�������5��Q������N�Kx�n.�F��-r��7��E8�/"�h;���E�ܵ�lyb�/I�o�B3�r�dn��6�GP�hp,y˩�PLAK��ΡT��[C�4��!`4g(߰�{P5U�+�~�&p�ӧD�F�e}�d�O��E3sNId�7;��O&rg�=rܸC�8%G�E�O�н<זU����)~���B�W\�!���be95�v��?���34��������j�U���/�6$�,JN_�vA�����2��'"c�	by�N��F	x>}$�0�Ӓ���G����y_�������|l�{&O�rM��A��
��AR36H �b�;X� _���SE���o��vWv�O2q�G1�sz�H�E�̂���cVDw(�݆|�G�6Z�+�u׿3:���O��ҥ����ۗ��B��~d��g���c)�TL�#
#�E�xh:��RS0D��~O�WؒTjwܬ�D	E}z��~-/E��8������J$"�?䀘@��8�K)��W��x󨡵u�_̚�fo~�C��W�O�b]Z�PFx�/ѵ#��i���e�~�[{�)��>|��I`�#ר�-Ă���O��6�,�U*����TL��\��FH��()
Vlo�nU��#%=*�]͵�?���uc�Ғh_?o��ِڛ�I5��W�|!a��$&�/�>�Mr��]W�D�KO�b�`�e�k�1G�t�ܰn�[	H�������$�>Ihǲ}�+�������r�Ӎ��}���
¿��@W��s/���N�͋a���x�N ��rįc����jNL���g1���cM悭�m	'��m�<�����Vk����y��O��Q��`(bP�t�2��S���ޯ�rt���8��^��r]�#4���-�OI0(0�e�/���S:LAM]B���Zآ#����HW�2S|\���]+�����y�?-^�+�\X�6!�,d�
�U�=*Mb�Š_?:WjKS�TjWF��wꕒo�N,3u�����HhyE�.�*ѽ�O10��4��6�cGN��V���iL?W�|U�&�2�����{��?�3��@眐��&��aL�O��J,��	�9Qi�6�3�B�9�s�.hz
��҅�V�Y�3PL/&�by)�φo�	�"�-@�C��}�Y�2�� Qd�B�
��A�EO*��=�Y��͟�,�p�A��mU�g%�Z^B��xf{��Po�#��e1�%3�o�K_�&�is�L��}O��hBW�`�Ҋ�n��ｴiғ+�N�=�K��/i���{\�#�O:��՛�74E���5���p������!n�d�J�c{A��m�լƎ�&��^� &���fƢ�|L�jK�i�����I,S�@]R0�	-9�p�)��ڹ��j|���~��γ�!�i��?!���NR/^l�k��a-m�iq}���%)�D\Z@�S�<[��ĭ��U��^!�-�p7����]����18(�-�ц�%Y�4������#��է���o�=�s"�]��:eҰ��I��6a�ͩ�5|�����]��~���Aދ��q��xa��s����ϸ�2w�1"{N�=D�J=��=N�Q��:����7'˟�;�OB!�����2��:�]#h"�N�+�������;�����7��᎑�On�9�u&\�S�x}a��w�i���a! ,ۈ	`�|�I1������`��0�U`���V{��&���E>��o-�������&L_���ܮ"5.� �}����;�=Iւ�յ��� ��vB�pg�
�R[���F��O��۶�s@_�������m�Qo/�� c���h�H:Ie'
1��`\�h��T�nzL�H���\.*k\��Ƽ�I�g���nM��H�f/I�в���j��@^�H�(�39k��k������-��O ]�V?�}��Sp��mi��Vء/�4;�R��oL�{9�;Y�Ϸ�ԧ���}�s@��AM��#�4#�\;-�˃L��0pʒ�'_�d/(>t*z��N�E����W���y�j���'ˤG���,=Mcv�^8�_�e�����9[������^����m���S���7E��?e�<#�T��3P��E5�V�\�C���D����烕@V�nlI���*�Z�ޤ�%p]���t�)��¹�U��#@����-O�r/}���J$�e��!��e��,�����:Iп'����S��k�:ީ7��e�ʷ�Pc0P�o��e��>�&@=�b������Q�V6x^�ØP��v�>�����!�9{�
�v*2 ����?r�?W-\J�O��έ��Fܧ�G:�����I�͑�!�.����L���q�R�y��U�B����O
 a;��8c4�62�%���.�q��~B����)��s�[�R����`�^�2z��G3I��n��+�"Y�TS�ZI6��xb�mC����>���\��A���pp�N��#�[���� �]H���{���)�8�c��B�����!������VSa��g�#|ÞċQ���-�1���50���_�:��8�GLoj���GG�㿹%Z���i�l*���0s�#���`,`���$ݗ�ѯ���vh�,C�7x�D��:��%R8,YB��� �춤��0��aD�����_��<_1W/�i���N��gf܄\
�M�^�DD�C]Hmg�=4q�睓�n��6�ھ��=����ChoQᑻc��|�*J"H�e��ý�q
mt%{����~n�H�ST��+�K�[^���A��;U��{���v��(?��n\@���Zx6_�&Qez�/�!���{���W^
�9�"�PB�v�M����K�k6�u�*����w
���di��4�����M�[H� �E�=*߅oU"��V��I�
�����-
ԃD�&��KSx��ҵ� �����l���Fs��laf�{�'J�$~���_r�#uw~u�V��<�k��6b��v���OHO`Xxq�h���;傣=H5'��'�?�1ő5�؇�ieB���`���]�g���%;ǒ&z��{�ݥ��|M�{O|1Pd�25�����R	a<��Y�����m�������~�G�+��m��n0�3����ˋ{�m�Ŵ�uu��	���H�S��svX|[Hi!�t5��K>���:Mn\AD���e�P���,/���ݸ�ᨬ'Q�*DdIG��M��ǉ_AI'����DR��ޡhCdY��L�d���
\�>/��D�A�\�B��혠b�`��^�Z�H��/��+u~/e�j�E�xi�;LW&Wr�;���z�����J[I8%'bp����T���a��ᇞ���s�\<�Iִ�=���t���>�N���I��bJbP@����|�9	���$��/�����n��M����g�5�4s���N�_�g����[j�)^�z$C[� �}��&Q�$�Xk.�gN�����M!f��G�6�2љG����X�_�ݸ��жf5�u��A��Aj��}:�8�>No�������������W���$�����_f��^}�%�y�Gl(lc���u�c=��/��>��lhcÌ/jzd,��U?x��b�U��G��.�_@��N�(��Q�|[&���ǆ���S�5N����ER֖����&
$�m�/���s��D��3��B0oӦ���S��8n:�0�(s�%���?"��E�Ȣ��9F� �f��C۝���_a��v��f�r�a�_T��_��������c5ڊ����)��v�C�H\ʍ�qm&�����Q<���5F��u�4��L�6�m�I�&i�p�ƶmۚض�ƶm~m�o��9�s�f��ܽ���;6�\�(]�z�tQJ�O �����n�G�u�+�v��%Z���r��U|�Y9����UaE�5�|r�1�gw���c���'�dE	���z4%ŵ�9�~t�{��r%cw�C&�%P��kړ��������,�g�A&��7H�d����*u_��\�aI���	�S����ZV>��}���2?>�~.R1�H��-M�|=�"�Jk�:/U�.�;yj���5�g���<݁:��8��d�{Fe��%�,�>fۨSh��LĖ*��BW���m����y��Fca������A��Tm��[�X��[Z���<����'@H����X�$0厉�޼3����ܚ�jf~UI�y��������!*'�Oz���k��d=�8��q�*sԏ[.��E���i��ḅ_�Ѩ9�Sx��7�~��|�ߋ�(��n3�����&c��=�BG@����kmp��i�{�Ŗ�[��r���o|����ɻ��SI�0Å��Y��	��%W-QS�:0N{ҿ$'.�^Q��`9y����*xR$���窵���S�1/�@ .|a�U_w]�~f����~&��21�t*��t���n����.yp_�uƠ��h�I���"�b:�P���a�UZ����R���v�&�8f�-�u�.��5���,������a��e��v�u�ˡ�r�����uߒe���2�]__���]�hƟ�������w°*"��q9�P�]n>�`ȧ̺�4�Up{eN�KN�s����n���覼�|Y�&t=��m(�df���LQVL�	������@����a��iȘf֯v��y?��x���Hxŷf���A�����e,c1��-{rY�N��Uoo�?��6��{0�~&�y�/�|��S�-��c�o?��e��j�`|��o�;��b���=js��e`�ٔ2'^��[���	Z�R׷��f��͎�����n�w,�����vEdB��6�6y��9J�q>��x��>S�^C��Ɨ'�lM/-���Q�Ë��6�}攩H�ݱ߉��
��Z�(PV��������]�O�'[Ґ�̰#76���x��3��jFx3Ƿ'ԟ����M�7�2��5}�<M�k��ȼ�c�I��t8R�;���l ���ʨ��UYz�����oW��黵�����$g˭	�c);ͽO��N�<1{�,�N���iNy��B$cN�M�Z'���ؓ������#n�5r	�ʈ����"�jtUG�Xy����-4o�4`zǬy)�}$	�@�/���zvO2������F��6�O�����V���I,xk�tn|୶=NvHZ7�cs?�EZ.�Rv����-K�Αy�/�T�Ll���v�j��L�>檱��WUh��= (�"��x��f5�$�h@鮞#h޴�=x.9^iֻ�#A��pI"=Ƞ��!��b��*(�\�2Q-��X�L��26����h
��I{�i>��bΪ5��t��I>���UL��]�x��cb�h����o
m��'���O�a�bEni� L�:�fZ�z�=�%�́���{q����`$5��3�Rh,$�P��[����y�իh�0׾�;�yDd�~���I��ܒ<̳�x4mQ���12tl��XW��ȗ�͉�L\���N��h:<�Zl��n7�+����sT�y??Ր���?Q��ďNFG�p���i7z�az{{v$�@����g	8J�d����t�#�1�𦊪�s���?�k�$�Շ�]�P����g��˿�;K�p\ߘ?R)���B��ǂ����)C�h!��{<+�q�,�� �ޟ���_>�yѲ� ��ݨ�ƹIK�t^���N�<K�]w)�55������3u��OC<�c��zU�/u7r�ކ����+c(��W��M��X��t�rf���{b��y`�ᣳj�4��ֹ̠-��r�/7dh��r>v�+���F�?�	d�}�vXB�# ��{R��ZL/!��e˕�B�]����yj3��O�x|L�H�z�Q�~^i���|���i@��t:���jV!,��FGQ������|ő�� 7����k�q�FXq�,��X%����C�������oǬDc:�S�ee�(Z��1¿���)"��b�"8��A�?��a�?Y������NP�z8��Z+-և�w|S�ѭ(ѕVlJ��Jm�ד�ݰ����z�P���-)��p�6\� ��+�R�;��>����N�{'��L�N��ўL�D�J���� �=�X�O�{�^P�?q��-��'��DXl1��Y���Y��28�]9���8	�]�(ҧ���ޚg)׽�Y���2����hy��c�U����k���,�r�m4����i8=����⩮֒����C�8���ngb����}�AY��:rNu�%��R��@w����ٻ�k!|�"�Ta��B��`���g�����c�ꢘ7����k�^���<�:��A��`��Y�I�X�;u�f'��L+M	;�,�qd��K��/���^�[@G-i��;֒<<�y��-�%r�5�Q~3`�nDBd�sE��_�$L�i�).����O��[x.G�[��_v"?X��Ӫ��%�=�)�,؛���w+�=M�X���B�X[�`)�XQh(���`�%QL>M� ���g��3}�g�@�
�Ii6�I��\�Qg�T����VF������~�46�L9[k�.}���My��J�liP�C3���lvZ�c�>v�>�fQݟB��H����m/7i�q.ٴt.����y����Wx�)���`��'&���`|��^&���p�ǳc���dy̜�',y))E�Ò, {j� ļKګ�<��#qC!���|�#;���{'�,F-,ڸ��h��q���hQ)�mܻ\��zG|�K|�J
���Vy��ҵ���a\��(��d;�,}�\܍0�x9;	w0��x��a�c�s|���zk��5.�^�l��So8�$阽k5�D��3��[�3	:���)Cj��Z=[�z�e�Äʊ�k���k��F��;�_��P\��.����#uE$�ʹ���N����%������w4A�^�;@��4Uő3��\ǹ�Ć���u���M���غ:��&��<�|��r�3�[V7��yPc�CY�v��98���Hcq�;�\�0ixt]js�{�"�I���j����S��\�>�8^*sX���o��9�"�X�]� ���,���T�L�Tca�b�RzJwf�h��z(���Y�8��xT���?`.��9��ռΔ���?�x����JZB��h�zMq]֤�c��Q(�	U)K�$����g5�4�(vYx��d�z,�}���r刵�~�d�.Yx79�_u'?�_�K�*C�������CV$ё�'�����<�����MURSGs�x���2]c!����l>]k�=��Wo�.�n�i�.=������5j��":0�<NfM]i]qg�R9+.~�5���_A'D�+$+Br���<��b���O���2����r��$�5���Rj5�ᰔ=-nL~��X�V��!�\�ֆc�"��'k6b�7@,}�����E�FP  8PR�"���QU��lRޚ�	�1S�E���BO�>��U�`���6�J��w�[(g��m<���&����q�{�<$�Π���0�@6=���C %�)e$ʹQ�R\$�Հ�Ν��M�.y�T�mfV�"�z��j������?ǉ���鱺�j��h�j��r+�z�������V�n��R���e�c
�������+��C���`�ED��S��O�%���(g��"�
�앨���T��	B3�p;D�������+�__���C#�t���a![毂,�p�QͺclX\-�p+%{�z��~�HmMZ6��@�\�R+���m�6��d��[��'�R���iC)ѧU��o�̭{*_f����4�|�D�'�-�/ܤ7��"�@��Ҹ�-~|�:�����e�;���+f�*47���C\�"� ��)M5�u�c�WwH���-�go
�p�\NA�뎭�߆P��>4�){��O@�GJ#�XJvt�b.n�vuPb����쟭�t)8g<�T�
�7���N��_-J}�lg�����}�#��|RR�5j���^���+I);mBm@���7�Æ���0�h�ת�P���p%�Q�44ſI���S�L���%޵/P���0tϛ���^Wc��#qv��7i;�?$M?Ў�%6�[���P���2������i����	9��Eb�b\��^o@C6�҈��"��+cר=oE��D2��BG�5��9O����f��bQ���пj�N4�\ �f�6�'�D����*�5~�x~�JTSo?�X	*�42-.�K+6�����[d��w7ۀ��,�e#��f��z-�����Mt5���FF�M�9u���K+0��Bр�D6�r�!4�"(Fj��E�R�[6�@�v���f��k�l�K�ɗ:��-��X���b,}V.����h.Um�O�������F[����+~~���sau4�Ԭx��N�N�Os����U�f@�_q��	���`%��T	�1	��(��&eY�o[{�[Uhv��%ڄ����)@�G2�F3�,E��;���ߙ�~0E���Tye�tsq� ��
_���Cf|��L3J��F��5ݱ��bC����E(E�8%�~ͯ4yB�[�.E�K�O>q��Fիmn]t��Y��|�n���֎�s������4����C�'&?NR�4����#1�k��TjRE�>��Dj���9x����>�9/e�ɠQ�ڥ;���9��l=�?F�E���q!��p6��萏'(�ʭz>@`�I���k�%�II"^e�pz~5Q���o�4���q�6��f�F�ad)pۭ�m�v�Ox^lh6��ظl���U�֚ �WU�[;�C�����wfj�C�����7!G�$�Ew �?:�5�0�&3�(/D@�����%E�1w�POw�#5S-�_Y��0z@<e�4�i�N�㸧ǃw��uY+���\�NR�?�}�D�q�Xd�"ڌ1�&D���]%⣂�&�q�K�ab������]�u�`F�h��t�?����β|�~4B�/ؚ3�
�Tz~f�=�m�_:+���6!�n��.���!VQQ~�2�ƺ��Gζ����Ǎ��)�����Cs%���b�����������x��w���=U0n�t�w��6b��ETY����?-���>@텽�.U�0��;�e�}0$z9���]t�Z���q�9QS���$<�{�4o�O��g[>�Y��pGa3�z����J)d�a������<�A*2��k�#v�w����`�@�q�o����-?ϟ�]��N�-RH+x9��]�I�ӫ���V#�ߝ�+�7ǋ�Âں�bA'=M?�d��n\���dIt3��쩥��'MaN�зp���㶘П���9�{[�ا�~��2�'�"+���>�n,G5��F��n2��@�PK��Y�|�}�QQÅ�'Ɔ���D��Ld�t��P�O�s)�v��ʊ� �Qɶ�����i�-��9��]"�����F<�:3E��~���·��S#����6�x��\����0���q�j���z�k��Z�&�X����$���Ōۿv|��f;.'?���,~���Ǩ��R�WZ���L�I8sA���g�<�1��G^�������5�����&˰�cӇ_D����Q��Ƿ"�q/(�e�{u����!m��e#W�tg�=�"�^yw�{@���P >m�#��\������8��<g&�Da���6�I^���-_�-��Y���y��Q�a�┴� ק=�O!t��P�ì�'���%��ǋ����qt���a����a\&F�^;߾�,�_7?WF��c��o�I��*L*di��if3L�v���=:���W��|�&q����P?��F�vO�������W��B=Ŷ�{�aL��[�c��3&�=G�I��]�	����;p�I���M^�n>�z,tyZ8Og�!u�$��?��G�~G�w}�v��m:���qA�a��� ����9���qv�� �����0�Pt����Ts��������&�a�Ԡ���v�+�\�H������7��!<I��a��]�t�8�֑�mw�W���DM��c�-
����6s/���Ua+Bg!dB.:##O���ߴ���1?,�\ޞArKwd�Q�q	e�ҟaS�$���k�1!7����y~d~�񌉣�}�"n#�� Bz]{��LR���$6�q�`4�g��HMnB����H/Udx�\���O��4�8�򸋩��|�1֠��bL��.�m���1�`�:]�z	��ɰLe#��*�#m�o}�z�=��s�df&X-��2����O���'��6��H��m،"��.��c�}���5�Gʒ�=�f"�r�F�0�y��Ϥ�7��]'q����O��V3gJ�W1� ���?�7����D3���10
WTTLk��������R]�����U0Ks�s�D���3e$Ŋ]`�_���)|���_]��L��H`2Z����v<�h�b?�{�ra>R<����P5�cX�/ra&X�4欄=��"k�VG ��8ԓ#�]�M�ϙ;��d���3�&rq.��t:v�6ݏׯ����;���1<ܡ��L�y>�=�P�43�ݲ'��Bݹ���ǽ=���^�w�6W/دqҲh>��ﲤ}��3,^�������Z�F����Ň�<dL�ib������Z�G��Os���Q�.爂̕?�����[Α�L@}��j�S��ɢ�8!
��[�;�(��N����i��C��+;Ф��Y��򾅴)�gl���AM�F%F�q��_���㡴F<��&�6�T(:'`��M����"1s�:+�V۴/�#FS#�g�gsL��l�Su�"?�\��α���eEpFJ�Qb��J��R�3%C�Z���3o�#�֛�
�6P���E9sL��]�0d�8}�}<콳,
Ү��(ճ"��f�P��~��3�����a��N�N�`\���Y�]wN���ߪg�Y䴐��2]�`*�%�j������=�a;f���g��G�iD��=���<������Ƅ���O�)��l���FZ��3��zX"`���5���� _EXը��
q�'��~i�2StUX���A�`���n���UT��aL�"�������X������`����fx�x����iZH0����~bN{��/Gѧ���+�N�Z�s��)��q_�hj�!ڏ��D�MB�o�{���J/[�!�\�#�T+�6I�n����f�*�-�ߜ���q����.Z�	~�&қ����A+e�Z7��|sj>�����h�G�Dǯ-�npl�)..n�)�^�$�/�%h=#`�-����6�&��5$J�r�gԞ���ǂ�w��S���±6�;�i�����Ĝg��f�FAr+�0�l"s�J�ԥ�,�r}m�m52>���4>�L���\�W�4�'{}_�� ���*B�7����5�v&ۮѧDx{,�2Qw�N̯PG�"��B�������y���<ʹ��WH `kK����d=��Y�OH�,����GD�ܿ )p��񲮡��E�������K�N��:��jQ�n1�\���k�5�I�i�H�8�t��L�/<m����q;��5����[����V�����X/o�>t�.}?��o���i>�gY��9t&|dwiH�"	?�w�i��C�K��fw�F��g��)�E�۷�p5u].�/�w�n�;K=M~��͜O���ߴO��=8WV�{z����_=-�.����W�V�������IأO|z�_�~}~)�O;$�x���c���
M�~��ܱ��۷��RGq���I�۶I�{,����E��_� ;�"�No){���C��Z!�T/�V*���XE#����5��}>�wݡ��{�D-��,|� ��M��>��suAo���~r��`�v���o9�� �iZF;��L��e�� pϫ�㲪�$]'M�}�aJ��惙ǫ�;�0��Q5�gW��^��S���iqk���b例��T�����0L�c��0��WO��y���5�:�y;��uŪ��A\j�j�\
������7b��Z~�D_�G�����G���ͱX��{q3�"��~�L.U#�\f`���*|�x�䷩j�����l�3B^5�jh"������~
�{����:Coz�8m.���������ә ��1�¢�e]z�B��e0'(�X=��n�!1 vv8���<� ��P�Re��0�*W�<~\�Z��q���Ũo@[{NG��L�k ȷ��lsd��|0�܈g�d�],��9Ur^r�?^>��\k��ۄ:�K����%�~u��퀊�N}İ����p�کKw�"��[7-���n _jGA���uww$R9m�^��7��$3�iH��4��ٛMeK�9	�Fe��N��Z����A���/�eE�S\�bI˨��Y�,Dv!�5]� ��-���{��k�q���@������D����U�qP�=����s0*�'�n������q��랽��^o� x��8�~���m�l�I-����j�����0����������-ǥe��9�o!/��S�������L����,l=?�}��o3AS���U��� ����ȿ0�x��&S6��E����1pE�����e�xv�escr�Q�����H7D�a-�e\vd���Ϫd��}��5&����Zim��WX��f�⒉����V��D��T򩘜�OУoY$���� `�+��5	���w��^��[�z�E��{�O4�0+C{{g�� $�r?�u����#�8�A}NԒ�)���~�E����u� �
�� σ����3P�*�J�qԵD����ķ`�^1�-�w�6�� (x�e�t�l�%�O�F��QQ8��QE���b����0�ʙN���)���}����)	�C/�9Ã��Я���x����蜚=�7,�T���@�ͶE��с��3̛����,//�x�i�&�I?!��1V��+�4��-����IA�L���0�3�!^(kC��1�3*�$�z¾2T��i��k��L@��)��C��s+7��D�Ee� ��܌�jk�o�R��4�t�p��}˵�}��0rIt��'tW=�	L���Ӆ�}�e��*7�w�1)��E�������9wk8���:�٦�C�
om7P��lK�6��ʯ�1��5�\�'E��E����S^�^NA���V6�Z��<�&��]��	sP�/� �>��9(���N�ғ��S��>����o�+l^����q�'���`/:�?p&�vp��ee��#=:?�_��PyXÜ��>ݮ�dH��n$�D^��3�>�o���L^�@�8>�Je�yiQ�&:�ӊ��%H^!������������r���V�
��L�1�YU���9UEJJ�n`�ԁ���9e��(��E�El�E"1�e�0g�z��âJ;q+
�M��Ā�	��&�nS�ҦS��A!>?�@{w���f�<f*�a�D7�Ĩ�#��3d{�~L߬� ��7 iP�i�FFO��F[_�[O<�`��b;6ӫ�����ta����O	|1��UBYo���k2m�s��4��������ޓ�,v#uRt�!ggl=�yV6U�g�@��@N>��0�K����?�RK%@S�2�A��5�ʔ���Œ[�'�	�z-�9?)G8��8��vm�a\�q
9�E�'֋3?���;�c��!˳\<����2���Y^L͡��0`��+6�=X�ڴ/�7�����J,p�Q���#�r��(����dA3mdD�nIvB��<�]����6:S�����&�Җ�ÆWg�C�����(4���(�lR�-eF�j�ZHoH�Mo�)c!	1۷��YF��Ѯk�p��z�"����<\h���^�w�ɝj��5'��U�3/�|g� r@_���W��Mg����?�^�,c�Z���Ǳj2��7�l}���!���� �[�c���a�8�g�O`>��x$4�z4�q�h��B3������~mT�~�P���P\|����͚��v^n�����WA%�5�"�1�A�
��	Hx�������Q�#'��R����$�hQ��V�BX/Դ^���w�ú��v�eDcH�P{�@�c?#4�O@C��N ����A���V���5�|�B��HQ��a-�ԩ�J�s�#���D��6���DV	��n���%�(k��}�\�A�7�ks���G�ZG�t�P��V=�'�\|Ǔ��_e:M��ں��c 	���|���̥���.������@�PS�SG����S��z�q�=m�>UK�3�z������`P��J��H>��@�+��r:B�+��u�&R��)߈�{�B�'��J�k���9���n�ގ,%�$�u�rһe �}�/H���c�%B�x�eC�-�	����h�F��~���J7MJ�m˃ z����Ih��S���0~���In��������5�1		g�O���I�����"����	l��{�콕����\9�.sɒL`��r�'�JO�>�!m����-�R"�{ח?E��5�B�|l[^�G�q��>��!0�r�:B��"fme�ħx�`G,
+�c����<@��$�6`���++Sbm� �/�4�t��}�,�����P����!��Qפ׻�n��a�,2��O�v��c�ċQUזS8ĥ�j 8���t��^������*��$C�6*i�M{�kn9ްX�#�B�(�Lt�3$t��)���A�^8�Vˀ���4��[o����WY�-W�Wot��? �1jzWy�9���2i]O�n�iʕrJ�s��軮^��s<e\Ѹ6D�5�&���S㫠	� ,*���>��-��`?8-���6�� ~����#,n�$����/g`��!#pZ�2@m�%��u�32�-ˌ �ԏ�/Qhw�c	�#v�����'EW�
͆h�2G� ��;�h�����=X��C`�$����I
��Pj�V��YE(���K��n�����V��z�ܷ8�f�g���9$ډ�҅�q�oǣ�`(���It�����է(z���������_�c���w��g	�G�z��
q�����%�jy'��'�,F?*^�.ƞ������2GOഉ�۪�jO��$������gL�c�eH}rC8�w�B�5��T�������U�_��J���b�����Ut�G���?���j��z)oh��x����.�s(-t�'�D�饒��o�E?�WN/� �e�XQ��B��FQ�����(��r	O�O�wţ~�.0�����V���'g��MՎ�¯�<���kQk��aP���~�L_܀4��r����QwZ���i�ûe�p~��:vQn�wo�ѷ0HȨ(���v���0���=\�����	HS��� ���}�^�%�H|M�x-��:�U�����X��m�M9.��E��r�ʢ1R���vq��Qʰw����^1N��%aC��~�>��f���tw�pb?�]�ܬ�V������a�u%Q�:��_�֜�q��k��2�A -E�z����q��3t�"λ6�����܈�
]m��s�v31���w?	�2_��������~��}���'��F(ۮ#`���
U�m� �c,d�!��UG���2�-��IUk��������L�`����<��m�ג���q"��ٷ��N���*���č��7iP�W�Q^�= �E���:U0�8����։:�%����ő��6R5ԧ�Nn��~�ʃ]D�������JO��XD�̙�t,��<z��)��Y8ω���È��d�C����I�/�A�`Pp���[�7��DiC=T��G�fU\6�dF��"1o�@<*|����`�Q�p������8�P�s�����3"L��U�ۚ �>. u�]�(2(�K�I��	��#����f��g�&(�:���-�g]�R�^o�sEOg�����$e��+-���T8N�L4j���_���g�818�����	]��e��/;��&�}���*�%Q@$�>	sދ�u�c-eߟ?T��\�A�� ����w4G�J�x�#4jv�TW��>��+�����؞)	����Q��|�P�py�C���⏭=;hi���>��ou����`��M�����ǽp���-��%����$K�������T�����+���)0��ӤvaxH3�M�Mͤ��@R	��N�'�G�h�ە��(�xG��Zn�F�ګ��v�����2���;��O��0��¨��A�6�X~ޒm���o�9luV�l���I���*T�S�j����q����F�H�e~Gp߶)a�d�n53��
F��ti���Gwg��M��~�=�4�R|���B8n��g|�c�(&�����+�d�Ĺ�Fy���"�<��@�I��R0v.������:�zsR`��L�\�E�t��<�xg�q&`�_��� ��љ�?�q�0#��#�Q`m����#�1���1Zk*x�zw�,�c�s���K�
��0���:r�=�m��ߜ����#���f�K���ŢRw��sa&�rx�[c��<����S)kk�L�6
�ͼ�����\�
X��-W�[eZ����ؑ����Ɩ����̼��mSy�wre
F����@�@o��Dd�U� X���|�B�vr}�<YA.v0��Aּ�z��1��M���!hm����o�m���و�O�ܖNö����y�G��p g�N�3 �}�m�k���C��NO\��W�s�d'	���ߊV�
' 3�A�T�;�i?��l&�)(�0�d��ߢ�e_Bz:š:~;z����7lEZ������JO���K�/F��!p��e[��'�j=�B����b2���Ud/Zh|9�nӽ��c�E����s^�%y��t��]�J�L���V��T���'���{��3�^�g���%W|#u}DDKST1A�||�CQ>ĩ�}�|]��z(��<�.1Ē9�t:
�b���Z_�����Mg?�	Ǘ� �����1�����Hd�W[~x��SO}�.��$DCd�Ս�Q�!U�S��'����1����P0�%�6�()���"��LL� ��rG�@8�����\��z����� ���:Ê/�i)�T��1�N��1H@L�Q�F���,��s���s�D�b��u�h��U��NR)m��Ώ�������&����s7�;z�(�y��뾥M.z�^	q�?���cB&!�v*{C�;e�;��E�:�X��R����_��&�ݔi���[H4��n�,��&Y�f��8���&�:�
��I������`2
e�I��������s�#��c�0b��0]���*J�K��w��6a�,̆٦�Q�*�� �<�7�5��(��L<χyw|�A;����l/�D��E�9��eZ���m޾V��v���9����{6����QB�W)}ٝ�졷
sՑ�#;��E�d{I�:���n�}�&���)sHp��觳T@����X�����'H�<L�Vx�״N2�V�=ܳ�9ڧNX�g�O�5M�]`s���8Bi��#�\��O�x�GT�HG�4`ͧ�>��(S�4Zf^2$���)���2���]�h�s!y�%yX��|�ڿ�SU<�t��[�~�|V<<��h�|�x����<`5�}�~�;���~�����wT�pm�׫�sg�����}9���������`,�Z"�B޶2��lPx��l+�����_�>+��<���-' U��d�"�ɟ���ӳY������ �����cFNL�hg��mڮ$�a!��ó�m�"����[ȋ'~>U���ܻ�k`�`m9G�;-AL�-`a8����+{U�����}�4ėAמ�s��N��$J�?t�a��p�}��dO(�!r9=���W��Ӑ�p"C0��.�;�&���M)R?L�
]o'	-�~��m��>�@�(`-�0n����k���%T�YgZ�/4->A;���߂����t�^��} G(GmO�oԁk�N*�Л�R��ɾ;d�������Q�������p�I������)j�t��;}���j�f*f�e]���Y��9.�{3hzM߅� ��$r���G��{�hF����������	����j26u��tdJ-���z�����d&��ʰ���j��<�(2�!�/��͛Ǐ9�l.16��~��-��{$7��)���e'np��Y,9�S�����K�Z�j:��R���� ��zU�OFw��o=�"�G��+]�
�GV�`��^ �a�a-�}���I����Ko �nk8�i���!;A�H"���I�zA�#gӝVz�H�mMO��WۯFB����>�S�T��Q�H�C���8"�1@-��D>�M�;���U����;:���0��+�
�OYf+���/��1tMD�⋵��fv�sq��&�&rxQ���5M�����ઍ�M��\�7���=�4`�
��ד�3bg�	�L�Y�e�7���ogS<|�#clQ'�Į��/}Sb�޳��=i	��ȏ ���Gຎ��,'�꣪�-NPp*.�	��(̨�:��s���u#d �i'
�|��E��Oo���6�m�iEލp�i�.��OP*}�z:�V8���͐��wP� ��<8��'����hG@���eA���Fs��@mm��#2�%D�]D���׿��c�Uc��qJ ���x���.�x=�c�DA�����Ȉ���jj�4��F�9��W�h��O�ƣ�����~I2H��������0.S��ʅ�����V��U��0uV�ǩ=�ӆǯ�c�����^m�p����ٝ��O�_��r���㈼�D�^$��f�K�&]jj����=b 0��8�ý�h���ᰒS��Z�b�`�K\��0��wh�s�+)3`�'�)2h�����C��d}�xڃ]4��ׯ��A�v�!ae�|!�<����N��M;�m�ʨ H"5��SV�rB4a�l�D0q�I�h-����.S�!�d0�C�k�?$L�rT{}��7m
�&qs����Z� �"-d�w�����~�s��x���VC=@�h��RC�`��2�`y̹������{qКZ��B1��.��H�aň�*�Z����ʕu�VwUߛVJ���T0�2�X%�F瞸�e���q+���a�/�X�W����hX,|�,'���zE�a[���3�|�����"_SO����Q�ҟq�7�f���>�3���ʶێHYG����,����A<y�^j2f|h�����t͍j��;�36�%�Ί��p�����"��㶘wg��5'�/���YV��H��HNӬgf	���~k�N}�|ڍ�]�|��H^�n` �v��xӕ���0�h�Ѥ������M�7�|Y���Z�R�Ń���K�Ӓ#�2����-��ڮ+H�a�g���el�F�����brt�ԗ�TD���'3��֮K�-3��M�W�ʉ���5��?@��ɗ%s��?K4���4���ү1u_���MH�Qp�R;6�Fd���;��?��hƎ'�W�[�s��3�^���E�1��� p�E������J՛�is����K�N�T��퇈>��0�;g���0{��l�2�J���w�?���]׹���K���]�;F�+YĪ�a4�p��Yʢz1��I�ar����á�!��5z��ڶ��&f�gZ&"���f��͂�� W��jD�}1�@��n�P/1$&����"�θ�@����'�
?�@�찦��ӿ%�X�����N.�
)��#��CՇ�d;�z["�����f�S�<�F��0}�����M�/���f�&3T_t2�Y'�A��[0T9Y���0��a�L�N���,��v�փ����:�C#����4@�gq�&H7wdđ����s�|�'	�)�H�K՘"�7����]2�?���&��q���ϻ�.�'�$�Be�MrW��Ϭ[���Q����@R̖�� V���ϲ��r��Ά,
 ���+q�i��	�F;����f3�k)�[��W�U!���%q�P(>�����k���	�N���Ipwww\��{pwww�d�%�{oի��fj�^����uWw��� SeK�&�7�7#��(o�&Y�O�|�?�Oz- �Wpp���.\k���[����#r�ڭˊ�>�]Lh�ev1P�����a�$89aܳ�7%{�=��}`2��*�	���%�yH�o�K�12�L����؉>������NRs�m8�ʺ���:'?3o���a/��P	󏖱$�o]�E�a2VO"�2d�M(j+�nkk���VT^ZBO���]Y���QTVVk��"�;`Css�AA�ri\��%b�^Nj���m��<�u	���j8��[�g����]���M�W`��vf�*$Y�c�͝���&uT��$_TM�(��u�R�\҄�P��|��Qb�5V.��C��b����:�GM�R̈�ӭ��
;��rؔ/��0�	>�e��r�f�D<�8�&fT�������SRR|��I�$0B�6��ě6���[f�e�,h�_n�wD��R�{�R�j���h��JS5ߋv��T|>>Rϳ
{��p�nH	�P�YZ�璪�)!��`�j��⸈�wh��d~�b,�	ۥ�c����3^�&�Ph�ya����6��]����Jk�%Z�� r�	��u�\b���әq���9���a��E�ߧh��#��wm?��d���*c�6:UX��N�J.�U�|���b6�ӸI}�Cr�1GS=,��G<��X{���~g�W�g��)��%�g�p���J��8�q>�M���4@�q�&��X�$������e�.�sIӆ��gi�o�ʥ�7��ܨ���������R,��t�W�!���{F���֤��)�g�������Q�5RGW��������:�$��pl%������J�i����/}����q�3\�fҩ~?#f��[�s���;�4�(��!�K�����e���*z�<�ZYWuff�)��S��՝�����l32�E�ڹ�4����tyvK�����;�_L�����7�bo{n,��}��NF��>�;Pu6����F{G�b���a��PiȩV��&Ưp�_n{s���xLރ�l,C���P��M���8�55g�q��@޷�'g~�;����>}�#_�݆]!��W��S��G���Q��B+s���^�3I���eFؿ:�kxN*�{��A-*c"�1�i�L��L�2���Iy�L�E�F��n+%z�*6�݉O��;�����{�����*��zaB@�+��`Z�rc�A�7B�SwC�>?�1)���\�rS��Ͼ�ρ�\�ư�I1��s�ʏ�\]kcf��>o��7%U�j���+�O��<�h��Bγ^��=�[�˶���V�/a��p��D��,3��Dx���Ri�k���C�MW3v�s*���� �L=� �i���s��բ���	j��*	~ā�t�� ��6���e�^=���e�WT�Z�Ao����r'#�ذ\�{ i��i��1Z�}N����T�7�C��Ge6��5�@�r��s�ԆR�m��� �ϤxP��b+�j������e}����um�I���g}Y�p-�|�UA�U�%�&e�$ɶ���v_[�<��˩� ہe�n��S����k��_��{��J���s���+ o���ɹi$yC��M{	��
$GQ����_���%qw/a�n�9 �&|��8X��S}��E�Ԩ���؈��X�e]_�i�n�v�]��K�"
�0�=�gğ�����^1"W����տ
r�ahNs���*��X6$�z������������ٯ83��x��5'�U]05��C�sv	����:=
*Ҷ(�8#���kM�]��j���IS?���@
EOn +��BP�p��?��jLGg��"�Ж�*�6wܞ��	mi��TesT�B;�h�������a&�/�̇/
8��h�B	VQ7䏷-��1�/5�]�,�բ����k��k+*+�-:�����i�.8���Ia��#L�ڞ|��_�CHM ��o�˿� ��b���0#�c��B��Wz7P��%-�?+Q$��" ��� 1>�p���n~gKY�0ɀ�1ʋ���T)�L%
���)Y�ӌ�u���d ~lu�c'g��5�U��tb��-����*�2K���������l4��e�~�7v���RB_���´+U�}3;x��Mud�M@����X�Ru�U��|?�4������Ε(���a�\�#���U�� X2����"�^��4QC���	��\(<����}��sN5���c����U���-������CȩG�#��P��u@�c���W�gM�Ea���V�~4]釼�\ [�4��N�I��/*���L�4y�Mb�猧��(���j0�3;Z��n���E2�e�86��8�/��*|��C�vF�U܇�υ�֩@3,ڭ�2��)b9��,��,��	��[�V��޲�)� c���=�DF��$M��fv9����;p��a�g@O����������kD���Y�5�͵B{C)����lgi�}��*Ɩ����K!+E�|��l��jnrn_�{i��ep����w�BME��/�NF8IJ���ةe�b����������/Ҥ}.*G�"�U�v��1���b�Śv��?^.�������w�j������������o������q]�͞c5�j�����J���xp��0�?��~�z%���"�A7&L�&�Q��ܻ�����w����`@��ۮL��4L�?"��43��0s>D�η��A��#O�G��_�� s>����Ѧt���A+��oL(J����o���[s����$u���L�K:M�Ī�����S���Q�H�U����?�?"�c6��T4�=K*&~��G���'��K���'��+�f�uUS&�R1-C�}` �(� ��+ ��S�U�c;|�oqC̺���#��ƻ�J���!F�:2����)�;���k��B?�3���ʢ�p_�*J���?���&Ϙ�(�ǔ��v�m��B�`*g�^��̐ǖ(5C1,�9K�#~��\��Y���K��D���Y~��IU�!�>WÖLG̈����Q����=8��W�f�Yu��7�Yov����K�j6����)���^�.m�	Q���Id���x��-�ӥ`\�0>0fRM��Wc
���Uu�� ��R�Al��)�S'%")��UWF�L��~'�6�~fA��8�r�W��3*��Y��Ӗw�oC��aQ�6�"U�]z��f���]�^��R��ً�����c��#@��ur���_�Qr���Ph���uƠ��$O�Z��� �ED(�����6`�KH'X�5�(L͉D���v�����r�@�k)([��{���O����#��-nc��0�#�)��(3]��%7X�X���o�Nɷ)a��������_��"R������uE3>g �b��U�5lĸ�W:
�s�T9�O�S�B��ƾl�U��i�s�P
�p��sd1&��qZnY�{��@唟�ie�h�Y~��!�d*�M��[u�P#�$�Jd��P�#��L(ӹ\�z&�!&��M�{^c��r��� ��8ؔ�ڂ��*6$���:���j갹�(]���H���WI�����_>����P������ov*86�4.|/<c�J�c
5\t]��P�e�Aa��BF�1�EN���.��R�x�88��[X)����HϿ�%�rά�,)�[��+�c1+ҿ~-�mw�K�Əf��"��[m*��uu���z��GR>��)�~G.�d�(46sZ%���g? ���cW�)�D�ܣ�o/q�{�>��� |A�Oj��-�ޣ� WV��d��K�D4)���_�w|6�3~��,���&���1\�r�̼�X�=�W1PgS���Y��l;���=˻W��*:�ug7M)���V�m�s���$l�|zs��>�mJpi�|���[������&��_:�|k��E�,�k>�N�5��?�	�h��� }O&����$]9�f�RZ�j3�D�46��j�E��>�9��kY>�d��d�"�%�OʢW���Xv���c�<�n����k/w�/��`R��|����E��h�m!ن��C�'�eӲ�-+b��L?<SZo~��m6yiK�������:���%�Zo��s������nH�����6pP"VrmfF�ފ���1���1p�w�H�@Ui�ܘjѠ��E�Z+�XBo=��>�'kNI}�8q�M�Ƴ� ������"'�&��S�5�jy��u���C�R6�AI�d�]�~���V�Y	�/�f	���Q�����c���`k�$gni�y���^F�U�Z��m���>��l�,�oB!GS_�������"P�������^.��j[�b�cc�"�Wj���b��S��o.�I�L�a?�7�HZ��䦃��V�eMm[��TvǴ�o��r�R.K�����|5�)���x���Fh`(����V��%ƭ)4��-��F@7_4[��:vf��C��-�6� ذd��ۄj��3��5a��䏌��%�)hmlk���-ܒ��w)��������Sk>
��*���2�%�Y�E�����5��u�N�_�y����}�d��Z:>���hyuu��aI�ݲ��(y�&ߟj���E.�+N���H^�a�X�-]�Q�0g:[�j*m�7Q�͸��+Z'Nٯ�M/e�2����#x����ʧC>��C�zS{�ݪ�n�0Y+ka{Y~��5B���9�a�U$���6^��=�ӟƠ1�����R 2=�?!>D�N�C*�6(�o �`/�"n�遼��-e��D��`����a]b�T�����;�������P����w�.�_�yKij�@��܋<����Ri���EW��{��I.���gk~��M-��|�AŎۈ1��ef^5��	�����X��Vb\��R��d�C�S�w��!�=����G�n��PЂZQs����]��lP�F ;���$nHI^�Ѽx[Vn�W<`r�~�$���R*S���Cp׫����F��kۖ_`!�c��f�7����i��n<��y%�D+64���b5a�)����Q�C�y�B�֫�9���������so��?��b��{ ���}}!��<gĤδ:Y�[ˎ�|}b�v�0�kQ[;���.v���g�M1�ߩ\;��E�<��)^��i|6���'���U?2����-���g�/up(X���Ґŋi�|��,ތ/B�IZu��H��C"�SK�ݻ��Pu�^�
��vV�2��+����*kLd�}?� �8:~~��0Ǵl�������?Q��umΕu켮��a�O����D�u��R1z欩��T����Kf>��}�U�N�sRzZ�E�fךZ;��d���Y8����j��!��� ��:d���nW0?��]v��Q^�s$�X�h[�����|E�h F��*����s�x�=�#�0x~��8}c����^Q Yz���:!UF��u�)Om����=�|Z�!Y�i�/M���"9]�)K�ʺs���护/J@[� ���I�&�s��H�L��6�P����:�KUqe�@�y��cXQ��(.���o�\a`��vWG}l)0��u�6���(��:U�����yQQR�='�[+�ߗ��.1xX�[b���2x펍a:Y��>f�&�6l;d��RC�b�"�1��p�}�D�9�q&k�<v�`N�8�?L�7���:gtt����VH9�����y�Rݶ�+�ۉ��=�H��t��?x�T���,�����W�6\d̂é�PE]��",��GJ�������u*b�ǈ��qdq�,�u������d�����5�x�v��-�@�4�/�n�ۇ�:��ss��O�g�#�s3���JٰQ�נ��y�%�P��;�7��A���5Y�g-e�n|A:ϵ�e�;��E�7�)�J��a��ۋH�6�#k)��KΰKz�`�1l��r�QN���oU���p\A��?��4���~g������/x_��# ��[��~�sw�BI?����"H>��r>SO7d��>�y�(� �,>�eY�4�s8����J��	zf?��A�,������C�P����Ǒ"=�;��\qoX���E�g��Z����Be����w�q���g��lB0���}�$������o}�<S?��1�`:�#D����a�ht_2G=���m����f���ORШ�%c�V/5A��P��춟R�ju.�9�4�.#�9�O;��6`�Q��Y��ό���v&��6�z�E�ZH�ᅦ�KNSO� �T ��O�[s����Z����/,W֮ax���F/�qϏ�rH�����x�dU{7Q�a]9��m+���<M=��<��3%J@r�<$�>��L'7�.w,:6�u�E���mD�ɱ�5�ߞNa i�	"[�����C��+�=`@�"��t��XYR������߫��-Vԑ����I����c��0�Bȏ��hYȂ�v��]D�2.�OaO��}5&U��=�w��J��%3,|�E૧���F��eؔ[� H�.ʊ��/�/w��*���G��e�hA.OZ\� ���;)+4��/���t��R�go�4��gn��k��_��:8W�s�9@*%X'H�|�[�׵I�E��Q�i|A����7~���۰� ��>|~i)m ���чt�@ȯ����n��|��U`߼/����L����0�K��9mVy��.��`�}�RKER�d��츳��KDۼ=�;4#�"C\��NGSt���O.��Y��������|�Y�S�S�9��`yπ3��a�����f�M0x8b���\��;ax6EMEETּ��헝�o��g�#H�-&�#<C�_���׿wm���dX�f�APD����<?�֖E��ȴ�$���['²�R��߫?��	�2��Br7����t��g��@kq��q�GO���>�����e�.Hoϧ>>/�-K/iD!*��x��{����m�0�v��&J�:�b�q_����6R��\IV�3�q
�-7�%���n�]$6�ܷ���<c6L4���`YH�@g�_JX�0=�c�T!����ݍ�c�c=T���N���<q�D�>��9.��H�� � ~�%�6>��0�n�((�r�^�߷���c��Tj�fo!aʜt,��F�=z7��d��;�8�{3z)Ρ������(������=���'�چ$������o
<K�}��U4���qX�Tw�|<��v�!�#Zg>�E/���Hy�=$|r��K���v��Fb��.@�J|�Ms�s�BO��-[�c�k�!mi�I��5*��mX|�KX�F��s)t����fx�q8͗�T��:�4�̥�r^ee��V_�,b|�c+���S�!����y��q���z��K�C�~��:�\�9���K�Q�v��L�a��� m�5Y���w��Sf�w�K9#�������U7�;>Q�%�Ԕ�m��A�^|ђ���T�}�C�
�`���oOH1]Q]__���0�k#��`���6�_\��i�C�/�w�.c���83ߒV�G=�������%��fȁ�f�l??Q
�y"f�����ݧ���3	N����\*|��W��N؉ ���bvLzz9����_�ǐb�nX��G��w�y����ԭ���o˺,���k�%����ʓ�j�qZ�ёS`�1�
XX=:�v�H{.�2Ja�V?Xi���kV�9ò�kUԠz�[��ݴj;V\��U�6غF���7��k�(�6Y��=�n<��T-����Bo!N���A�M�r�U�
�/a>n�������I8����������y�w7W?���)\P��:v2�B�?:�:�p���I�q�0�u|���fQ�:�|����"�n`��Ƌ�o��^�+/(\-D:�_oeu0�֒:"H��w\&E&�ein��Y۹WA�?Y�dҬ��3y�!���4MN�d{������Gv��B]�HLÊ;�SV.=���8������w���~���m��&�P�K�r�$�c�i.��UG�g��`���sۼT�_%��ݾf�#��p=�r��ǖ�/�¹���
%cv��z�����2qܛ�$�몤b�A�K�����[�������6�6L��D1���O��TKl�j#��;�j`���<7+,�zV(�L�N���i���U�.�z*z�|N����xI���sX�g��Nx�=�w�h�R��-v�.�#��i�U�}0����^�a
xN�?gJh�HN�|��s�8�t{���+�DaV! ���)D��0��+!�=��BYX  ��w�i�"a ��qw <C�D����Vm���8b� ӯ�K]����k�-��8��4}���!	zx�s��'ڍ�w�]Z׫$]-F�w7$��q��m�]?���c�;�7�1��R������'|Xz�Q�S�����d�#`���K�T�.o	#�_��e�+OR�z��;`3���vT��L�o���k���\���nF?[�-��N�Ĵ�ȧ�L�-l��V5���yh�H���J7{my7:�q	��I�sf(\�b 9Ot�f�W;�`��gn
���T��z{hyv��(h���ވ%����O��L�8��2�J\HH( r��O���/������]��u�p2������^t�8l8l'�q��Zz$$d'���B��4/ƺ��.A�Rc�5s�L��L�����9�Ԇ�qbs��q}�P�qߧ�8}f��R��1�y��y�m�D����:�%��^ �W�JC׼�v����MTbM���Y��kT5�f�����]޼��o3�2�-��Gե�{�Vк�m�$O��]���M�R\�r��68�+;Dw� �&����iv\�����ʂ�@���\Ϸ�C���AR����>�yﯖ���͇����?\)O� ¨�q�N9��km
$��sh1*CgId������7}#���ϑ��&ֿS;�v��"U8#�Ƙ���B��`!)zw��D���E�D����X��������g��H�ֲ���QaP����f2��zB`�M��;k��6q:;��X2�*���[�9 ������NA��������&���c�@�I�ͣ.i25�)JߙV}��|��Hh�|�����۾Ȗ�#-knld?n$���I������%��;B����f�c�l�\��2k�o����I����<��v�f�=țy�Qi�d���=�0s@�,Z�w���YL �4)���yO���𝎫!.4�wJ_#k��
��AK�t�h��rV��[WL����3%�6or�9�q�ц���m��C���%#Tī�ڗ��6*�G�_������}GO���Ʈ��1hV�:z�%�
�6~[�t��������1��J�vq++3�(��n�.]ne�Z��.Jy2���_9p�e�q�7�E�����v�Ds���͒��+t��\Yp(A��F	"�F�^k ,;�>�_	�M�F���|g	�1��-ѻ���"Z�Lv�M���\�Y����yB���� ��,o|�M��,��5Ң��L	����{Q�]#���<��!HP���A*gt���K£�|�� �+��u�5��x���?n�&��K��[#�q�Ҕ����h�)��BoBD��A�3<��f��i�K�4L
 ��U��
xT�����a��Z��/:aY��=�w�>ta�<�&��w�~6(4K�I��k�/Tx����y�z���<�_�uq��;W��46��=�kyVnM�6u��Vm��w>?�~��ūU��_�w7���R�̚N�`X��%lv���GdR�����L��^LVZB���?v�������-�B��ۙ>�m<e�tY��fm(���W��Z1Q6 �0�S-�?��{!��X�0��M��#螑���~����(�[���00��vkJ͐���8A����Q�6u�u��-sxr/m�ǚ}Y�i�H�eY���(4�Dk�y�K���v��%��2�3��z(i�c�KV.<�r&�m�JpZ�<,k��'�o<���'U������ȡ�M��������'yA�B�]$p������t��|�^��U����6�f1�<? ��z�	6)ǃ��D!ӌ�\r��V2��PAU����g%��PW�`t���CD��-IA"��$����"�4'�k��#Z���ٺ�鴉þ@����v#�^�%�H}}�q"2X���`�8��ַ	8zy?�HET~N��gK`�g�����l�qDCs���m�p�>�H�����E�|�{�#����&��I��AW��8�,���8���Y�[ˈ�P=03�y�}ḗYGYs�R�&J���O���f������H�1h�Y/^��.�0�Q�Ob��i�¯Ƴ��	�����j��U�@�$J=�pr��Za��DW��/(��y11�ppO�-���FF$�������� N���L w�YgW�w�b����y&ۜ}�&��$n	�V�]����`���P�h��wB�[�
��D-�����9>G\�癇0k�r���2����N+�d�#��S���د^�Ƚ�77�
Ќ0
9��0	+FDI��ժ��ͣ�>��4�l�%�D��s/��Tp_�v�|%�.Z�q�!����L�s�?j~\�v4f��C�U䞐�$��oF�]q�ǉ5H]\�	ƹ����:�X{��M�	\P`^�,A�(�n�#өcuh�m:�Gh���[4�V����-2<u来�W�3�>8����� 4��^�X�f���jU���|k;�\w���|~��&0
�\ل�X��!�3CE��(��C4�_�?�d�����n��D�u�-�թ��⅄t]Eת��d��>��J>�jTY��!\�\�w�fo�`-�^|�k��ݱ��`�	 ��:+,�(��5�C��
 �BLa-���u	C �R�|By�#:[q�J�P����Q|	��b^�!,��S��Π�c�� �du���)�c �/놷�loG��m/�,6�"�oQ���S��x��QE�� #��E,K�W����φ�"wk$`�	3��̅�xtA��C�Z��:<�YmĐx���I�?��$�_m#Z<Ϩ�	z���*xZ׌�J4J�s�s����)�V䚞�6�`�j�ڧ��E���,�%�o|Oc�#��S�/mABvsR>�����G����C���'���3��鈒MF�r	䡂�A�PO=(E;��ߣǒ3;��A���YP��̊�%�|���э��!�i{Qw =*�6E6-��(�,�
J�|c��6 ^�E9]����@�� ���"���5�؜��[W����hLP�����$�!%�c7I"0TLad^C�Y��%Ke�7���'�cˡ5{����^�Nk������?"?/^�X�bXad�k����a�������2o�������7�-������(�-�b�cL���QzX=�q��w�$q��\{9#����*��S�R��)��Ї!�H���r���I�S��q��/S|/����.�cq�p��r���< �d�o�&�L��(X�[N �PI���ʧ�z�w8�@�O�1���M����K�v�D���_����O����|p`A�c��c��m�qG!�`	ﴋ(��KS�&�	mF���
�5@�H	���0y��q��
l�MI=I�)�$/�>m
��6��c�!å��������ԑ;|��8��(�����ٿ9�;��ؼ����W�*PW'����4I���d�4 +2?;d�V�$C�nSx蔲�K�\�;�=�x����k�`:��MR���ᚇ�s�3Y����x���4#@��v��&��drSx<���.���(�}/Q$��}2��ܒ��8������Dd��1�z�v�`�|�����3�(��(`�;w2�+��CO�h08(����WD�T��0�i�]L����.�@Y��E�-�Z�n�<�)4�J���̼~)U�W,2�i- l��t�c�K�͍e�<��w�, Z�w��+/]��}oo@ ك���9G�����}�G�,��uϝ���O ���;���vd˼�R��#r�ӎ���4 �bkPD�i�9 :>y��w���h��'�H4Ҙ	�|�%��1�z�z�渽'��dB�9���_�,�L�O��6�����vu�#��A�#p����ÄAPUM��#<��
A"��@�J���:ݡ\�ti��̞�h-<�P��/f��9P�]>����7a�eO�v�򅷗'"b�Ԥp�Q��81�w�7i��j��Sʍr�'-X�B�����Z�Y���W/������Y��+�f�����v��jS����&V��c�؂�����enf�5J��Ӆ�`'�����QQ|�h�|�K��Vɀ�ߨ
��`�a��8�� �kHN꣠t��ϵ �)�ȖZт����� g����Jc�^�mƝ7��a�=?H���0� 9�v���{q7������Ktxˀ@:g�4��Y�!ÙQk���mˆGVnDl|Y^�H�G�B@ ��@M�7�����g%ő�aT\%����0/��1#P�j�,�h���aY,�@^�� �d���voU��N5���Q_�EC5�jГ����_��t�I��L\�T�Y��Ŭ(НrP\0������w9��3J� �(&�W��#�)��Pz����A�sr��)h�%�i�IhG��T��F �,D����m	zfB��ih8��z�����3W��u�}�¯�.��?�Ev[�:��j�B��B�/ɪ�o���ܓ� )7�Ȑ��I5`k�,k�}��L� I���hQ�Z������p⎪%Ii��Icq���{�E�y3׭����r��%��돜G�:`�0��gF+އ��5���(���c/��L����C��fGi�W"�N��O����"a��`�й�}�̊t�"! ��e%D�.��� ��M.c}�C0v9�Na��q��0��X�1Q�C��o��1ȏn����m����U-�Ѭ�V������X�CNPO�c7�n'�)bZvx�0pŎt�W��� W�Fk��&�� ���e�߽x��P���ԾC�?ņ)C������������C@CO�?]��dk&�ω,4�#����/�)��]���ډMFݑ��]#���7��/�/�qE�,>��(�L?p�Y���-o�$Gz��q�bk�� 1'���7�
e�H��g�HLo�f�5�zg?8¤Db�zf�	��yX�KZ�ao<�T���^.X-2����%�>���Ɉ��C���f���rFJz�[`3>�⥂�K>�:����)Թ�s�.D�V�Ej2��`�@H���
��Z,�u=Ht��~�z�iB��!��Gq"��x�f^��/��x�wt�9�X���4��(xx<qWгWs��=�<?�Tw��f��#��)�]�K��nJ@��mީ��ȫq$�=D�g���UwU߽��$< �$l .,<b������=�
L$���l	�	�`Ɩ 7�
E���wK|���hۉ�Q=!Z:�vӇZ���E�W��_9�-��M�����'�$)E�]���#�Ķ���Γ2�뛐J�[���Plk�Z�
d�C��	F k�#H^�� _ &ܣҤm}~��pa��e�%��=d����9)��[��U�1���?6�6A����iR����B��.�G�QR�޻��'=�1�m'4'�\c�����L����s�P+2��j�޻N����T�{��XaF�`Z������ ���Pi��軩�)����u�3.�-�H�
��(�cHC&%F�6�KEO ��b�=��������"�!���x�4
A��F�S`S>�9{e1j���z���t_���!�[�z��N�H�����F#2:=Q2g�zi<@Y�C<�e��!Dr�zG/j�<�3 ���J0o#��Hϑ(yv
/�p�h�q�bi�b�@�v	��!��UI�ޱ�ށ���i��媰��׵L;��R�����"��F󳇏�B`��r8!��+���'��5p"�@�B�-L W��6�+чXQ8e��q��~�}.�c2�\**��^tTk1��B2#x������j�Fd�ˁE�0�x�q���Dr�1e�e9L�fkw:⠃L��� ���/�Z������,�4���l�Z���
w\{C���]/�o��RX�0��D���r��%��!����`���$�"0]��]"�����;0�����ǐc��a�dS�a���_��:�P�NKF�v����B����x�S����<���S?H�N�`�B��LR��E��)�2��������5�!�#��,}�@ ��B��"Kdw���%I�4OP� <�����_x�c�u�qɵo�Tr���艹Az�z`�r����'D���%�xP��+X��\�`Q��2M
�Wm/�-LA�����MK�s�(�bEn�^kU�`.� )�B��|*o,P�a��곛XRH{B��7�)"�� �C��j��2-n�\�o�FT#\�2�������Vý�m��[�B�aTS���<�<�7B"�?��/S0�����,[%8�����C&,D.��;�Cǽ���N?�2�7�������橏�\!��HO
W��k��o���a�?����|;�3>�mAz����i�|�睥����B�}����S3�׃�!3Sr0��}�>����12�F"8��~A�Q�G*0����#�F6�c�Ͻ���N%F΃Ӈ��H
�;~�]y��{b��]Jf5'P[�R������6b�p[dpu�.�s����w��V�X�v޲Ŷ�v��V_��	��`iQ�F��g�6��s��؎� ,�{N���c|���̅�e��C�c����ؿu�c�����k{&t�M[j�+�a3�ν�y��9���w��p���A�$�j�f�*�=*��{�����*�ƭX~'V�I?Wli1�
����|����=�"�ٞ���L��~��9�����Ң�,����ID�ꋼ�ۋQ��cˑr6���<=BIl�)3�Q��*�����IZ�#Ä��U��պCU���qTK�X�(hBs�;������K��D�������Ws1�'u�)c)L�w7${�}�r�j���	�Åӡ�Wr�1���Vr���t������dŷӇ�kQ%��+U3����8�F���%^�I�g�}!��כn�Mݚ��G�p۬}u�^�.�c`D1����Ԣ�LMj�4@
�>'�'��[.kJDU
��w����	4xe+]� �LSp��z`TZ}"or݇M�����v@��(�)~���xq/VZ�ٷ[|ÓD�[�a���NM��C$���h`�5� �����&#w��a������H�m21}��Ua����~�9*�{�>8�8����ϴ�"�UD��#�Ȟ�$V�.�@��Q��zhdL�D� C�+���E����؉J12ɍJ���m��<	>����g�C��f/3ϙ�$P�8�ߌ<+�]�@w(EJ(�������	��}X�#�F2	n����b5&��4�ON)�A�p��r���,43�P�_	ʁ�c�@N��61G�I��[���h�Ͽ�v=օ��\|A�
cW<���8x<�z�:�싂��]��^|��(���Ʊ>������v%P5'�(58� EaR���P��٠iz�M|$bM�[���f�L� �{#��|�]Z��,�?�'��)J;;��.,�f�G��;3k��_��|^�'�t`�+�eE��|�̓,2uu�D���.�L@yCa���P�"N�&=�_��~Wz��|^�TIu	�bF�O���i�H�!F}g�?�$^���~��n�������id�J�oY��Y�0�f��>}�q�j��R)�)׿t���[�_��	���w�}�JWKs����N�5�a!�q&
F���N�S�	o�t�}�%(��*~�^���K*:�d.,K�?�-��{��~��XM����;J<JD`�`�䙟�,誶���[���I\YTvZv(@`�'���Fd��Wf�u��7 ����0Wwnڠ(N��Fg�3*�'+R�}�l��L��zL�Yv�51W���O9sO�=q�j��t!�����RuY)�����4[$R��2�XZ-���wL*����[����^Bua��~(֚���Mȹ��-��b>��UYQ�*F�>2�Ee�*�m�������G@����"�w�:g�=�](a=���,z���cta-���UIso�p�W'���\�i��R���h$�AC�cr
�)�4jz���Ź�����Sks����M��Y�jÝ���\1����j����W��=_Cq����ݵ�P�P܂w���P�ww��n��{y>��޵�C��;g�왻w֜XTU(�i�O�B8�״�W���2����8�֝��oў��ցa��W��T
���Ⱥ5��
���S��0��xOnx�QD��8�&����&YHc�Fz��{vI�)��ƺ��<�Ds\P�,�e8�b��bp�����+`�_�V#l����ب�&Rt��<�e#����J4��P����fS�@2^gW�H:�!�7U^N��r�$���o�a������kT�~&WK{��)��Äo��{M_~�cp��\�p~H��t/��Z�j���wdN�.s(�]$�?_4��fqQH�ٴ����m�;�~(���Vw��t��n�IE�Z@���6ύ%��[�/�
=d��4���]�7c:�hP�2rU�rZ��)�P��z��C�����|ԣH8v� <�4_���rS:�-���b�x�#�v՜�|/ɓ�7���g&[��݄�:dE���q�:x_��4B�R���_������&Ku�
������Vԁ���^�?Y��Ӯ�xmV��ֹ�o�'s�>����hQ��'��r	r6Jy�-ͯF�y�{�Z�)�����b�����)�)qt�>�Ϻ&�q봞g��~q+,��^����n�D��? ��X��$��� x�(��Y~���%,	���$Re!]�9��"�oj��Τ��>��z�$�C��XC�]חL�V�u��D�����gWX=�k&�wR0�4����*����rL���r �J췽�o�԰ x�sE��ZOg}���� 4��/�R�ǅ�`�I�V��Gw�E�|(�ct�>��#�{O�?�(:a핿=�im�� A��y�g�����r��[��u¦���8g�.>�1UY�)~��ǧ&{�mM��DH�L��s�QH��{*g����<�1:Z��)�$�r�%:@&��k,K�$zr͆ņ� ��@vMj�I�pC��̗�Le��?��2����mm87�@{tcgd���������8YZP��4Y��_�﫵�Ԑ�9\T�w��UD�^v�uƖ�F̨vt�WC �
���U?�;y?�E_��3���sͨOg�5:�JR[*7@���dx/�E�*���KE��-�m$��C���24{K9o�C�@��R��	N�f7�X�Z���Д����zQU�#��tn]�8夥k|���+?~�ɦ��G|��%����S'�<]���]S�h9:���&cQO-1H9aM�l�鸪D*�����a�M�2��8��	��1���?幸d:�#�dn}!��#�X�N!�BY|��z�|Fk��Ui��=+q��b)h���;�@����(���vZǌj���N���s���~�,����s�����	��1��f�!b9��4qX�g\\��Ly�b2��>y~���f��vc�XC;&s����==������&�R�jf�<[��+���w0�T��8n��"���e�����t�Cä�s�m�C��!���/E�-HF�_�8���o,�02%;yt�=��E�2/Ezvɲ+~��ܞc`ċ�p�P*����en�1e �L�� �
Ɉf�I�1��H㿺�� ��;e���t����b���Q��4�t��+xmn������~�����/�
0���*�\g�Ѹ�.dum8W�P�-����q����r�����*�^,���`��hm��k�B�s�K��^���իW�#չ�g��M3ZU��5]_�Q o��SefC	i�hM���PT�]T�Y��y(T�_���l�i荁�1w/�>�@�8����Z��+��9�#X]��db�)�ie��t\�àL-�(3��(=7���bZ��O�m;� !���1�r(g�Ǹ�#-���&�����(X6�1�:6D��D�En���|�J�G�6����9d�2�mC�7s��*!�����b��?!���(#{�n_-�v~I.:�L�$��>N�_X��1°�_`��=��P8��M�9Ӝ�s��,�6�8w���!EڛfldVν����7��a�,��|��[k��lJ�0����	��R?�?��E�L��~"�p����m�l�d[�������#f�;M�N:�\0�i���\����վ��¾�0v�V#�u)���&.���T"�B�b��z�]3���4�>��[� �Ȼk"f�*83�����޶S��
��^������ŀ��:iYu��l`�U/�& �|�`I% �qC�/Ac���K�>�c/!�
@)[������H
�ta/��1��X��S����*��Ҳ l�D�v��,v����|�d��h����_�c��/����}q���1��څ���Y���7!�yl%en�a,.��s �UΓoͲ��2�*�@�����"L��8��� ��/������( DW�B��E���P��F���+���.��Q�IzS���uZ�C�?& W���{x� ��6�z��ˢ�7��=�˂'⣸��)S�Ay �$�İ	�B���*Dc�|r���w��}��|�Vy�gA�d��?g�U�(�1�)�ŉ�T�76��}�lN��3oM���OTUE��(�(��A�C��fzu�D
,�c�+y����ͺ�/x��Mˈ�����c�p"��B�����  ��2(��9��%Re�v�R�9��H��7(k�HKh�f�N��(z�q� �7��$/����U�3G"���O�OC��&+C�{8���� �ӱ4H󌛔R��4��M��ɣ+�t��A�2�1�>3�L5�y7#����d RCUE����0�ȗ �� �:�~X)x��8	L�p�}E� ���=�R����T^*^31<A"��~G0��nX|L|Pm�| �q �1T�wn��`���xZ�J��,�u0,���kv�G�a��"�@F���x������BV	L5�6����0��p�
S�tA��m
�����抔V!�a@���܉�ɺ����s�Kv�@	�4�cß��B������
�{�
���1)��&�(���.��E͆ /��$�f���'Qg)ݪHcCȡ��<�%�6�*�S&L���9G���7��J8|%6�������/�)���y�%E���r��yH���PPTE��Z�[)����l�9>���D�����3y�T�'Q*��{��'������o�e�9�﯂A�6�:�1)��<	�`CL��l3U�?�=��ʸ�t&�r�x=V4̐�^p�'��'�/5�V߁DJM�e-�8C����G��Ĥ���/b%Zt�{Y�b��~:	E
�%����x=�fr��~��G.��(�Ai.���.3Eo��sA[���(��S�Q�(n\�JE�R13g�H� X��p���|)E*�v�ˮ��M��C��Ā;���X<h�q7�2�:�:�+ - �������01ajg�w�̤V՛o-o����ѳ�#!^�v�o<'�.s���+�7�4xi�>fJ��1*�{���°�� �����,ZT)ѓ����LdW@?��ٙT<>MAsY8h������	ɰ6�4�sn��H���\�* 1��O�Eu!n���&���06�q����f*2R�!��?Hߚt3p�?�j�h�MFa~�"��F�אd���"�����5�����[������K�%� (7�P��0�|�HHLLf%W $x�|JH��K���6[`�6�p��@_B��#�q�1�i��OV������O���*��1&k;$5�� ]om0+��+�{�h�r�Ϣ(M՚'3 ���d0��U!�CBuAht�CS��}Hx�������B���4���_U����A�+�DKΌ���p�$�7T�)2�ɀ�,�������H�|�9�W{?;9��h.5�����4��9yE���q�����z/3�w3�P�.��f���Z]9^1�cMyI0�H��j�p�3�.���ﰸb�`���F���YDR"I����z����E ���}���*LF -r�&EA��_}bx��?��>?�O1\:��YY�y�8��,��P�{�.Y�Hw}�ǇU�|Tjz�}cy|�(�6+h�����8Nk.~�s��R{e]�H0Z����Y��$I8K=�Ua�u5��7TQ���%<����a={ךS������t�gM�b�bS_��d���
ƫS�-}}:�J.�����Ɂۋ��o�VGA�5������[V���d0�5��4-?����SH[9@�r>��-���m�2�b`s(F�Z�m��!���F��e�^~�����zu��$�`sD��F��7��D�l9���}{C�{��������-�P��{�ٍu�+B�������S��/g.J��6)Q�ү���N�s��g���>��݉�a|W�t7��>��6O��������/�X�h�jLN��]�RL�%�#�f��x�^��'��gE�9M�eRg�8o�߻H/H�h{p5XB!��0�� �\r�c��P���SG���%k���n��+wH���[��%`Ž	��c1R���E�W���Q�F�����]�e�I� |{�o��a���e.�vG,+:슦_��|KV[3��j�%h�?�����A�7��Nq/d�LѻL��-���r��©�+F͍��6�QG`�=�᎙��<G��^-�>�O|�������[h�?�L�L!�!�*�$h5=L@� ��ϕ sz�D�'����/�3�:�����Y��(ߓ~�b���i��c���&H^�sH�|Z��E���怯��.{W�E�&Uف�����y�ߡ\+�[�&��l�l/Ks�{�ץ�N���l5�B�����)�����L=��(�1�Øa������6]�:u���GN�ݤ^�p��nW
_�6��4/�~S��QN��O�h�7ή1r��n?]8���w����3E��l���ӊ� �֍h	QM=�a����ԉ�}qF���c6��J����s�)����\�z���]p���n4l�4֜&�PI��Ķ�	�y��I�-�+׮�=��/Tַz<�V�^˖�=��9��lf�a{�w:E��@�1�N1:}v��mN⻿|���{]Js�m�bd��h��E^~�h��E��k��9�Zd�.������A1��.1f�3�"ia���3ۅ#�y[�"(`G؇�n<��g�g�No�m��`�I��#"mN�~mmǎt�e`o��TOl�Ŗ�*��f�$:�Hү�f��=��/?�=��L�L��}�~���
;́�3��xo*�s�I���cw1&�?�R�c�ŌS�k`
1���Vb�������-S�J�s�hhi�)i���D�kIr`T�?�z}���l���L�����c�/W*g��WG!r�5Y.�6[!���PNB�#���i�k �H�.��8�_wv��1I�/��1�� 4mAh�*��GӬ2P�Z9����xj��������uy؟j���9�t�1�򙛼�q��o��e�z�|�8Q�ީ��BkR� ��rD��i�q��q
C )Ծ05~EW'�%"о���N��߭�rH��|ׄ��l�̴Pb83PW&ђ#P|��$���C��<.1_#)N�-~��i��l�΅�����H��à�U�8v,3y�յ�!����z�q���,�������$���O��<�|Bmp;�q�`���W����M�<�v�G���0�j��Cp\�`�N�@2���$Y�����V��-P��3タ�U�����s�\p�1���E��>�h�o)��'O���-�,h�AE��TX�(���K�mА���Ņ�aN	���6�-":�2��WfL5�p�.�4-8~0�@�؀���)��#J�Z���@�z��Q|�\����)(ʡ��TS}%�d;����	\,����0�+�"s%�����p�/�������.q�R��=�V���[����H��Ѿ�ݥ	IR�
���2��B��O	�K��N$��^P��X�hU�8���:�F��O���3�!�Hp��ط�k����ef��@s��r�6��f0��;�L��~*#6��j\�:��kJ��i?��8��V�Pt�?�y7Q�ﶮ���"ؔ.~�e�k�O�潩���wqڊLT�̪P��ⴞ��0 "VAbBo����L%��r���O�ǻ��q6s�P������AΚ6M����u&��&u�C�}mp�DG[�巪�HEDʻpX�"0L�I/��V��P��qM�)�o�?-iȸ;9��pP�}� �
I���o���"-�6�Ƭ�D|�u?q����,�cQ6� ^m+�Xa�K���U�YG�@팤P#��T ���ь��O yX`�v�	�T�'�`���n� �vf���e����D��h�d���ݞ!�{�f��/\w_�Ո͡2�_'��fJ�r;��tm[�D���?X�����b�����a���5$�,̤�Yg��l�A�ղQ�b^8����@�2؍�)/k>���c�$�<,\\�/Z�sߟ/�Ff�m��*iH����$�\l�"4CO���Ź`<$����j�da7�V�bx_ia]H�џ�)�mβ�m+OU��o��ZO\qƔ��OQ�{X5�'h�G��0�͐iS�	P���X>%=�sT�P�9�&��0�Eî6ͣ@R\daW�}.A3`�w�%�O
��J1a������֪ x�$x�7��%�Ka����]��h��F/:f��|Ƣ`�E�~�S<qJ�å0�W#�#�QbCDU�r�zw��+&k�p\�DLF��Y/�Z��G�sSL��P*v��#�[d-�r���P�2�)P#��j-��w��J�3�~ů���`��� �4���_��4�Vz/��i���p𚎠�%o?Tcz��h�>kE��@M|��q���f�L�H%fH�Q���(^�?jI��L([l���`�:䔩���;E/��	�����^QQ��E^`z� �k��O
��?�����T�L�'��A�)�'v�3�i߅��b�T\$U���{�� ����rDF������ʩ��L��xp�p�җ��@�-�j�nL�6˂�|�'*�q{�5@d��n0�49���~I��%4r'5�#S ΟW��� \��a��4���7�E��F�CR<�-^�+jU�# �j~N�_�,g5.y�C��m���t���Ӹ�ŽG�;2S������$G����a�����#-�)닟d��\!��eG��A���ZI�c��(�-=���;�rv��#�Ǻ��Y�`#��~B����F4�5�&�5�&Th孹���.5_.�2qZdBuT���W��!cJҿs#kk��/�'H�u�jH��:�j���S���FсDG�� }kY����J�=m��Y�vd[:���d�珖u'Hh!�5f)K|5>䖈"%.��%�%2��@Hy��Q �n?�N���o"|Ka�\��{��&0�%�#R����DqE}����T=�p8��5��Hn=
�7[��emA����k�/�ҨFĦ\���r_1*�4l�+�s���0�[C b�	�ѭ�*��A�-�R�K�*� a<���B��6w���I��-|�p��WmQm>��4ΰ��Xǵ��&���>0%��8�՞��{)�`e��`�F��b���\[�Oeqĕ�)��H{���d�����S��s0M�p��9�7Q�q�vĀ�Jw���H��9"+#.������s�Db��R���+�Ɲ�P�*��L��!�帶g>��!<,������C��ڿ`��\���̅���������L�f�/�Vvr�@o|�_>��󒛿ʚ��X����r�{5{7P��]�$L:ŝ�$��_�I'X�Nj��6��A&9EReexɘ�^'ѽ�Xs��^v�p�.��ݾ��Y)�ʜK��\z7WȀ�^~�����׉V�6���V"���İ	ؑ�xྭ����	���������v��,��)��P�Op�b맧�9#OPD�y"��@CLXƱ��W;�O%�G�K'�[l�}�5��tCٮr���R5��T��i;K�-E�˿����^�e�����ך�!��Z�gGխ�b�t3�x��2ݭ�-X��'��]RP!����rK� ��|�b����*�Z��w3/��{��������#!�AM�/�	�֖xY	����պ����]A<�x&#O��̹ڻx^��ׂ�"���)�>\	���Y�]�硥�&�&j7�������#�!��S�+���:�|�� ��'�U��wo���)�"ߗ�s՟�y��S��i�Z���bv�n-��H��tŜ0^�)�lqF�x:.��T�=��P��z����ΐ�����kZ��`�����=n�2����<�1�k�ż��hg>ҥq�u(�5��vEI�
_.�lo�A�h�m8���2����[�gL�䣝�:��w�*�J~\�Jr���\�tn�`k�o#��G�T��EFo ?�no��'�� \���9��9�y$dg�zŌĴߝ㉋O�d��3�E�f�;s0�=s\X>mG/��#�0�U89����U���芤��^�pn�	�E�!�	{����9J�S����Ɯ�٣�MO�`0�� �aR8�N���9]��IL�ZW��䛎�(*a�F�'`N���=���ٍ���h<!��/�����;��,���\�U6�ɉm�C�!���2^�_�}�P���<��%Edۦ��^@��n�g'@[ȍդ�zQ��Y��ž���ضs�Y�1w-+.T�F���V�߇���'痄|�B��.W<�nN���e�U��w��&^��\���$5����}�O3��b������
�M�rrý�E;;O�Y����I���Cb��[7M=c\X9-�@�H�.�q�h`��Zs�!���t�/���P濫����c���/��;�a�$����Z�#(.�5�@l�HL����?�P'JJ�[^ڈpח�%x�����~!�͏�y9h|7.���w�|��n��o��҄i�a�~�q���K���a�|=�8�K6JtL�ϒ)z���$��d���T��t�� �[E񍍔Z`)eo-!l�`���rX%Ӡ�G���n�*�,�n��-Da�D��K.�Uޝ#>�eod�kGҶ��`�M��z��9fN*����W�Zz��~.�*���*q4�m�U�#cα)<6������Ȇ@�Qs%V7�������݃'�����N֓8�H����t����p.f{� ���Y�H&��Mv}�r�D̮ל{�%�hB�������O��vM�ڈ���\`��ݗo�����'|�p�|0���D�/DԠN�s0�l�E�Rݘc��nj+�; 1ui�"݂�����g��a�%�bᚤX�����/�9��hr�U5��N�s�ΌY*�a��4k.K�a3=���p���d�c0�M�c� D#��LO���ۿ4��~�|�,M�$���~��=�Z��?����Ф�O�ಛ}���*� �6sY�3 �Z��X�=e=���1�[���# X��ї��&���f��ld㖤���E�c&���w-�3��0����X�M�)���R�w��#��w�� �2�#���=]Y�e����GԜ#��$�����+R��T�v6����N�R{O9�(]���^{њ��F<Ҟ'�I/�3��j�i�9O�Q��{��YEʄ;07zVJ���U�&Ɨ�U�9q��ɣ�i�����i~_��
� �bEt؂����15���C�w�h�����Q�"D��u�3��m���reI�k6�8��QV?�U���������(ٳQ
�5�M���j�d��E7:!Z��QD��Ӈ�b#E=7:8 f̓u�?*��e��x��X���I��.;0n9���\{{R�]�鎍�Ш���DEn���rR���O��0od�&4�b���i�&D��}F��!8�7/�%z8�K;^S��S<�0��n?~��$��[����)���as�H���ϗo�\+
أZa���z#�ʁҨ���j����ֽ����ځ�1q�6��^��\�!1��rs����ȹ��9XG[��'�_�6S]�%	���;��θ�+�B��?�;� j��!\g$�/vdF_�N�ګ��3[�^��0����C�,K�K>�[�*��r|(8�5`b�jxby�>�2.F�.e�Ғ{9ۙ݊��u׊o�z�����{sv1���Fi�:��nx9��?��ȷO�`Їޫ4mm_m#�YuİFk��Fڮ(�\|Ww�����̀�������_�6,����i��"�
s=�!�8��r,�A����M�~p�c�ȗ���A����Z�\z�t5��o��>s���cW����4Il�cW�ݭ�ܧ^�&�O�;�~˕T�w�Ea �Q4�#���%���@�-���jT��Pr�)i(��E;�`��������ށ�[�!1y_?��v"tY?ѝ���#�n	� ���m�KVB.\��<%����؛���v�?��kxW�_x�E�S��-�:U���j��az埻�}�������\�]y��(���I����厂b�|�q~^��k׾�����e�^�[(���@����*9(��;��T�ζ�ڳ������H� Z�����	{���KJ5�E�r�'.�z�v�tq�t���� ��Ȋ5�*�?�ƫs�9���Λ������Xg��G��y����j�lm���cQ��ԩq�UR�g�Ay�D���K�''{�͛v늺,���f�Ƙ��j���مYs�B{�=7#�^˲��	�mk�{�̍ݟ����(k��袄�F�����}wvF���jI����W*�$7ج﷢����Sn�~c�o�MULo��:>�I��DX=�����m+�!B�����v.�>�ƕ�ԧ�y=��E�BѥV?>��/1�����i��ζ@��=����Ei;Co�ݑ�	��~;?��a��\�PQ�;�_� �����]錘����|����Q���WX�0�f�5���Y �:]����ΰ�숸~�2��	�����V��r(��+�,�U�k�BYMl!o��KV�Ǆ.vW��O04�ҹ`�쀫Š���]b���m����"Ԇ#Q&�5��o�� +��UK��Ճ	A��,K8K>İ����6>i����=,]��_��ם��aDp��8Z=�j���-_�w,ޜ=j���.��|w�^�p��3 ��6���;<~W
�@j�m��h `�=Q�Teo��]}�s�Q���L�F���ѧ�%�:��-����:1t�H���X.�\
��G�Gw�f�5",��1�{�}}��Ζ�B����H_�/��ʑ�4�����xe�\7�X�J�1x�����(��5�1��ֈ?�����K�^">�_��ѷ)���2ˉ���;oBH���T���%�f�BJEm�w������cu���Lփ���P�!4�sH��MO�+ݿ>0,��\wgGbĿe�m�;�N&��c�;su�*�@��}�;׻�SSř^�b��>�����[���Qe����?>���؂/٤�Ηp��G�`�9��
ԅdt�ܜ8v?�'��h,���S���n
8��zmS�`��d��[z]�|{֧���F_ef��9Q7�$�ȉL�KO�tz���O���}��D"�e��r|e=T�ڰ;7\��7�6FB�/��L�u)R��(s~�bk~e}y��_�(�~���ا�k�s�h+�L�)��9ei��ɠ<��^��&�O�p�T9�4����֩�����q����ohm/������R���nz#�%G�V,ܘ:�v_"z �@�1�����9��
L�����j�����d���"~ ��`��%aE=��p��Z�s�w��õ�m�x�n��퓏;�����٫���F:��B(�ئ�����IB�����`!#��F�s��{�~��ؑ
%*lHK]��yUb���"��J�Q+ƴ���vO%0��z��&��hD�	 ��D![m��;�-�G9�>T�]��&Zl�(��o�nY���7縩�`�|/A��"l�ХU�"���(F����B�¤�K�7�N���@���vH�*]Pw�+�η�E�@���i.��CGwT��^ǧ���|1aD�O��-rΊ��g�+�<�r���p���UȮ �Ӂ���ۥ�	�y��o���8͟^n���{��kgG-��ڕUod�=����i���&���!�4��uI��U���.�C��DH�\��<7�c�v�P���ABr�DǚĚ�W�S�0�)+�b�6���쏞�/'�njG!�f ^�E��^!/:�I(�x���<1ؙ�s�2Qfu1��"�����:���n����9�i^��G����zb�69$u�X'_���T��Fҋ/�]]dr�6-��XɈs/Fw�{���4��I������	lC��#<�ro{��r�nwg��j�9�l�mP�RsD�l�����O�-�ڃ�:�ƍ��M�^�+;{`��mDW�JDԓ&_���%��F��Z������.����{�#��Ğ�w���Qu����^�gZ 4NS�7L�
K6��e����u��]aڻ�!vZ&|㼷���BtG�l��$GnUQ��0Sh�Ar/�͟ywP����n�.kW6ͮ�P��&VA����_�(���?�{�k?�T���@ʦ�B���;ew޴�u��!�ӰVf�4�G�+}^�L����Îf}��ޒ$B��������]D�AE1�6����t�K܇����C�i���m�n/Q�r^�r�&�"��D���_��E��ڎ�jt�{��V�!2q��z�V�*Q�F����o�>I��曗�<�}�2�T�M'�#%:?�إg�2��M�h�]r1�=,v�aΝ��ګ�{�Sa��7u��.?�%�����։4kN�T�&�|N�B�<2&nM��)�o����K @�ZM��o)�ӫ�y�i�C4ߚz�	m��F�M蟺ð�Ǻdh�!��.�Y)/��k��L6��2�^�Yԡ�6�5��]1�Q��h���l��r�:�vW��#;W�J�mɌ.���,��k����P��[��[d7����c��=�`��8����rUV��aa����#��D�b�'хJ��a�	�u������|.ƪkݑ�$�~CFq�W:��Ee��3	�i���Z}0�bQ���̨mj�/~�j�u�c�!��7/J�C:d��/B�)U��y�L/����*��\D>���@�9�l^�U��`=��`q��=آ��/�p�DjM�=��xl��bF��*�	:j�/ᶡl�d�,��%��{_v-���8�L�D���T	#+Y`!��v�w�4f���Sjf���d���8� ۊ��~�XĭwoCA@�(f��)�h�es����`���|�`�@2ϼr�A�(�Ҙ�v�]=IDuvy�|i�|�=��_�
�5��+�5"�M����c}�:��tx%sۀ)1e	�+d�3�I�
�b5�"���6O|u-�5�\P7H���zA�|3E��Iۅn=�'
��~oE���eŌf&����e��$�p�s�|�Mr�va���in�����k�r�#�'�4����K�#=v�]�yk�og�Չ_ �^VO�o�C�O�t2F���ڗT譿fw��\:�s�z���k�2G�ϥ�D���q^-/_^I�srq�P4�~�g�� Zt+�v	ҿ�|2 �N�v]��պ�{!�N�q{#�\xi,d�$�%b�x��m�ĝ`�Y�Ux�=��j��j��	�&fBBɠõf5w>pţ��8;�{�Щj�tH�x�qwl uG![�7�s�h�/��S�8t��-���j�d�"��Թ[@����/�*�`*�P�n��������e��I��#����;s�P�Ԋ��e�n�n2���j��s��d$�[�..��vA�"�5@Jf�8�����f��0�-(c�OO��-�a;�����]�j�Y�cw��%G���X�a��,0�a���T<�_V-���|�b��"���
�w$8�s!Qp�.��r�U�J�e'�݄"�tɓ?�j�M���zg*7��!��<`G��ڇ����L�	n����	��1���Ձ-4���?�N������+�� 1B��-0N�v�é����B,鄇��۪��X�}�nA]x�G�oz�z}nl[�bU�c�!�&�x8SC�ދw15�>�ܯ�zj}�	��f0!F����<����g��z$����#���^H�R1C9���}��Tw�Z��\`���P�)��y`j�V�/f����zk�Q������3��-?�=�2.)w�Q�Ϩ'_>1��&0V���h����`)�P�lg����׶«�Q}����`RpB���^dg7.�������'�1��>�h7�=�q���W�SG��7�N�ﳟl�C>;�nU�Fr�o�G6�}�٫�7)���s��&���e��MC�c�@��ꓻ�~�s��g��t��yB�����</uNkr�ʃ%/5�nb�7�Rr��˖O�U�rO��ן��P<�����6J�ns���Ì�+��r����?�_wA+;#��Ζ+oq�0�&v�瓧���|��wh�QA� a�f����W���}d	�_k��ϖ$6�-��N�"k�j�=5�5��uy�m޵o1��;KWA�g�
���v!W�-B���Ʋ&D��D6�:�?� 5��M$�:�Z�{3��%�ֆ�z�Ϻz��6-�z!k4'>�D����g�h���홺� ��=#2'�~]�ֻ��Z��"�S����	���].�����z�+����K�~���%�}�S�[��ȉ��!^G9Za�Г�1�-C).[$�P��pR�$��Q�j趵{鹉�0��F�d�v��F���{H��o��J�����Jh��+��FqCU:�5��]����f?m{�r�e��u�8@7��|�vY�F�M�[PZM	�C��T�,��O���������Q��_>�֤K�49�d��Ei�����yQc�����?�"��(ʾ��^�]z��F��3h}���;�9��!�b�r��6��6�
��&/����������l��0� Gq[976����p���a�[g������jn�5s��MQ�Od�?�a�Jի;��f�H����H�k����b4�H�31'uv�D���Y�䪳a̐
%؈yF�����`�%^�R��}��u�¬0�k�\���X�S�6щ^(K{��m���"�g���(2�� 4�ќ��HL���[� ��d��w�O��h`��0�"C^�M�o�q���~b������bD�y �&���&T|-?���l�̢��O�O3���0��w׻�g��&n`C*y9�cО	�R�T_i��h�<�:�xR�|Ƙ��]���lM<j��>�u!5�!d��p�i����Y��ӞE�ԩ^����Gz"���J�9'p#��4u����I ��M����a�����I����6�sW�)i9����ml�5g~�r�G"�ʺ�U��V���X�~��gp�tci+e8����U+��$�1�����������/�L��/&-mA���-��g�����2�'s�"W����H�+^�d㚒��&� �X:晔�'�&�f5�{2|�������$O�>,N���B�Do�S�Ӥ6���鋎�?!�fu�o�)�~��3��1������w����f��z�r�ϝ�����d���#��l�ci���Db��%�SS�V����;8#IV�f����D�}���"q���Wt��G���[c�"����Jj6g2�ɗ�s�D=�gJv�=}V1Я�6��������T��*���	R�ǚ�M�7�P3�\�����kg3 �Ydy�cfM�	#�~��NW�ۍ`�C6N������wbɵ1W�'�Y`	�ñ�y8���dH�j����q��@��&��j�n&-��C�(� .�:�F0�A*x��V��ۗ��� �4~��k�1�"� �b*U���ը�9K�YߟN�P�1�t�A[J��C��(muZ�]%�J�x�uy�?�X^������ܶ�T^���}��2��ȂQ��OV�����p,�N���O��X?^�� ŢZ�1h�FbR&�$ba=�[���vm�h��8��M_F�S�LI����0�F���:�lmK5�(hq.pL�T�#��5�R�
r�|�/�$�~�1�>�A�٩�E�B�r3����Z��!������l�?m)�n�^T	��օ�ڡ��qCL:t=Oi*�d�l�!�#7'�N�d#�!�R�_�����㦍K*������ܛz���5H�)��? �@^�0\�]�]	Y%pv�2�����+����b���wyν�8$_S8��x #,G�YgЙt�F��2F�R/;�7��ǯ��qx`����Pkm.�<��:{�#�*���[�b��e�^��y�
����I�og��'Dʗ�!��ϩ�]c0���>�n_������.v��s����w��w]g�\
��D�������߱F�q�~���/������|�K.���������
W1�J�R������cn�1�Ҋ��;O�Z�-[n64�����.X���8�V����P'�#Qcj9�o*|���X3s{�ݎ�,#�3^����%�F�;����^y"m�2���qf˛�w�����@F��
`@'�����=��꼥|gLjr�`~�1����p�G�9����.)�|n�y\�#!f���6�l�4X��ପay�!V�4r^�T-��8�M}�u��Y��H7�k�}h���XkZUP� �����B^F�\��B\�u��(�C6K\�sU3�`�k����%�A��^��m�x
��/q�>B����mQ�"gn�\8�z~Q}=\ ���2CnC��6�)=�?d�����e�>�����c��{��P�)Nl/N�B�;:�g�M�S1^��F�$�§��8��Ltl����VC�{5̒�yuV��e����N�֎S�#��j�WgU��m�ַ>�����p,a�f����j�(���DY9���-yh�h'��"G��<v�IZ�� �������ut��V��;�=�־}�A�n��	�s���aV��'���k��d�;�s6��h�j�9�L�E{���.�8���/.·��\:y<��ٚ0�72��������`8�^��u[������� l.H0\��2���\f�u�D�s��SȔ� O���'�"�/v�C�@����N(���B|�{/8��)��m���(Av�َ"xؿ	�BVy�3έ8��ˎ��?������Mk(�P�2O�m���Dڠ' �1�Լ셾����kxђ��f̠�]�Cu�\b�z�a<�n����<`&+���9���n��l��A�#�{� N��Z���qE��/Z��:��H�8C���1�Ⱦ�e�r���`���pl�+#��XВ�^��U�*O9T�p�O6�ǲ�B�CD$|�������׻���&g�g���+Ӡ�b�1d��!����/2�{:xd�I4Ԍ;f�͘˝�}̒�q�ӑ�0~֤�]���6f�|W9�����k���2E>I/�X��2B���~�}�<	��m�xέ;#�j1ؖrq���cnZ� >S�)����L6��g|>_������2�b� �HI��{1�����|S8c��Ʈ�A�.�����N�u�X=��<��a[��';�Z��Z�>Ω3ojM�Ӿ@�F;��k�t���٢�a`��Q%�豬���F�U'�a��'eit����̘�8�N��w��p��n���T;�`�����x�64�.��4/{r�^f�2c@�f���Q�C�pd�2Ȗ�oo����8�u�Cs���9�;��͑�+��u���ZD�f���>+b�e�>�g�t]������Y9�C�L��W��!��+��µ���?����/p䷵W�y������ʪ
�2Y��! 3\�2����N8)�<8�)&�玍&m}���h��^�"��;DB�Ce�k��M�r�[<���"
��UG%9f�ϛ�bvatG�zÅp���ls�I��0@R�{8��$��=�!�8|���p�{!tq�"1����a�J��A���5Ív���6�����ƌ��:o��y�x>�H6����vd�(�|�$ȞG�	�%$y\T~9�,^S���\��%6R?��0%$8�J	l�OН��j�"���=>f���?%"h�Q�Ѽ��w��B�V5�8���!��7�+G%&��mß�W@�!s�]0Ͻ ~]�s&�f��`7�d�m�9 �p�όpR��w�k���v��״�u5ǳJm��A�J�`�_D^|S�8VC�#�a߹;�����V�w�̽겣׌}2��%қ���7Ἶ]���~�{�.�y���3�4���7���awͣ0!��\�x�@#R`�59f�a��u���٥Pﮀ���)s~N�<�Z#�l�aFFd#���ƽ�>�q�CUv<�X�B<��*T0�⤊c��B�u\�2b�����)�@:��kQG��^b���.8Zta6~�p�s�}�Ie_�ࣖO-��h9��+�X!� ;�c�/�0�^�������=<��x�}[�`e�R�n��BD]{R�^���k}X�0N�X����̷�;�e��W��m1���	���c徙�� �/�h}�;F�\�w9��x����ZYvQ�epK�5p\���6��$��e�T��1��W|�o�)Z;��`vv�5�f\_��/��{�^쬄��  磊�S����^��f��<QtE�X�a�'�������((�Ρ�\�4>#z�{)\��W^��`!w�U�>\w:�U}2���K_l{��g �k��w�����ϷO�\sr�yP�����=��*�gJe�DvoK�1p��m�%�$��E��H��9�"#P3�:�K�酹Ba�t�O*��Cm˸[���8�"�0���[���������ß�®�=�@�kq�*ϙ�]�]����L���:/��$�|y��f�k�+�h�c�>��X���4�F|B���-���=oA	3�T�^H�����A����1u~#��a�2���=��w���(�8A�eϠ�`������pTY4r���=�߿�;��u(Yi���5�=У��t����_r$ϩ�$o��9�	�&@�n
1C��Fo,,���Lߝ�9X�,�T#���Cy�4u_��AY��_'Q7D:�}w���̷1�p���/X9H1�JW�6t�e�/"�n�HZ�F�C�A$Q8��bE��\��5�i�3���h��.���N[^�M����_��3,t���E��S�������`G���)�v1àVۣg�mt'˱� 湪b"`�pC�+�_�:R���TDTI�2BTg����ӑ��=�^���)�xιp^���������w�Y�?���y��Q7C̓�i��p�p%��o,��7��OB�G���Ȕz�O;��]�o�û�8*l��m���Y�������=��\�˪��yT7����#naxw����ʃ����z9��^W��a�Y����`mh< �ʄ��U���`͐_m��	W��8D��<f|�:�6|�YD}�|�&uV	�U���q�����YFS�b�r]�Qɲ��U2hu���(��Y%]�~��V�3`W�
7P̳��lo��fB1�Q�����)�Z���v�X���m_���؅���ƴyp n�s���A�}�k{N��f҃�M%z0QQ�PŔk|�o�-rg}oѥ<��q�"�!��w���c+���$���!8$[�%���!8�h!]�q@�S�?s�m}�`?3�VF�A!K�V���V���Y)c@$Rƪ����+�J�Qo�V�oK�t�\��d?&�V��)�eBl;��^�i��pPVG�E|�s��<ߝǍ�~Y�c���^�}0{���>�pOA\0���-��wv� �4�;�>��+	�25F���������sj������o�h^%��u���/XR,���R0����]��6W̠5dW����H�*e�zG<��_ȓ��Gk�59�ߕ�rg�>���?º�e1�ݸ�D�16�@;��6�Y&�*���)�[��y��k���*΂�JV�<6�#���<�ㆮ�pk�P�����Y
��Xg��ֿ1Cl�G+�E��;��}Ӿ���Q�*��P�����5l�ݎrh	t��>�R�̇F_�0��N!��}�x�	�C��*鮉r��N��mg�^��{� ;�.\G�qf���u��g`?|BF8+��({]̘y�M��|��>n`����Aw���l�jLeO�~p�Q�ڞ���t?�[����򲥅�B���7$f��轫���0bW��$�#�Sd0#�~��to��g�v|4Vt۽�g���^aH?�����	�C��pJ�0�qD����p̀�}����v����ٛ��|]�%��h��qfy�g+����F�s�{���b=���f��Ϟ�5�+y�O�\/����u��2ݪ�Cy��Z�kC/����y(n�]'�!���ƛҰ�]���}�°]����Ş�G}b ��=S*���w�
��in�:���g�a2�B�[��{��7���1��)���~�_�p2I@ֻ��Q������'*�����q-c �ލA�r�x����Ǡ�=_*����6�ή�����ۘ~;��ѷ��]��:�j��P�,�%�q]+��}2�������<T�UO.�䚬݃��6��x��4%��2ybu͆��8��ޝP�U��8���7.f���w�.�W�v���������;.�Ӿ�pG�C�{���s
g�0���^����,�|�|vO�٣��
&_���;��kp�R~4�ʭ�S�)�H��9}��M����^	���à\g*�}b��0��'�ux������ j��~��А[�=DT��׺߆�7�����yP����y߁�7�OU�s��l�3�/u�k�	��-^�e8�5���+wQ��5��j�;߾��p�Z�9<�e[X��w�����pR�����k�3�	�d�(1�@;�$2��1�2K�a��]���2�g���VC���e��A&�C]�v�J41ڹ�)�� O�J�b�������'`�K(�^��!f^���ٚ�o�ZF�mU�y��Y���H���Ⱥ�U2�N��3����ݿ�e�MQ�4U҅������A1��ڻWX!��8���x���+�B�p_�}7�3(fO�1�'�) �C�EYHLd�$s�r�����m?�΁n@��-]A��ҿ��������A���hf�U:�����oö׺D��$���j
#�����ؽ	Nt�C��r4q�0gPc�^5�ߛ0�)K?h�~�v/��\�g[nLxO�k�}JE���(`��;�w��Sv��v��@�R�x:���X��4`�i<�S��Ww��_�ɭs��ջG��{*p�)>X'���M��!�QYX�m�������c-���q�e\j���a���b��a��	���W�~�=�D~��3���k�$�~�eC��G�I�m�����
߻�n��e��եE*<"]|�jg�Y�ŹmJ]&���`��X�&]G�qWcDZ#s���;v�����̙��$�F��NH�#j�t�b&ӊ�1�!S���7�8g�/��	��|]SW�^
ˆ��?��?d��>U�V�ȱvіry��B�H䓼�!ܑ�m�32�<�
�����vcV��fg@����kAr'e���Ƕ?gܵ^��S�������sw�H�O�3��g�l�U�����/�����y�+!G a��󭐃@Wt�7�<	�]�P S��G|<WٖH'3xE�Zn�ES�D�c-��a���i���M˿�}��_���en�.ﮃ"f�uDD_�����B+ 	F�C��e������;ކ��5�ᵟ�͛0W/����G^49_�b;
����1�����i��H;�:A�p&˝�*7]%;1J����������L
�[$�EbL9m:�Ć�Ϭ��?4���(R����ƌ���0��2���o�4�|R�W3qy�s]Ì��F���`S�띥��Q"_w�|8se��Rn�|Va�T&�{\cU,ϥ:@�vI�������\+�{D��.o���c��h���=�5*���,w�e���O�q�E�(k�B��{�ѺT]t�:������Sƌ8��q��s�@�4Fp���u|��8�f��0��/�l�W<R~�t��2�LYa1������d�JH1�ؙ�q�E�*��<:,���=<@l�Ȱ��x�$�8rb����c���)����LI�\{������T��(6������۲�)u�27FF�{0��S��YE#���2}VԵE��0�E�>�U�ߴ�s�/�eJ׮#K��oZ/{��˲��e��}��ȫ�2�	���C��8��ױ�du���w		�^��8SX�*�	!�k(c��Iwq�$N�5C�b��u���w�%���wM��Β9�:�s�=oJ���Q�ېg��f���H�
eP�1 ;�u�eL6��%���sU��=(٨�I�o�����Nb}��6s z�L��r�P�5u��^<w��M�X��7��V�,d�|���%�߷b�σ��'b{��̖�8g�>v�������Ы�-��%��G��ԻC񳒥��J^c[?�$�/X�����x h��R��x���Z����켛�s����e�
fD�d{w���\y��3��!,�_��?}r�C��h8��88�(�۱��ɓ��C�.(��g���L��3����S�@C�8-�ze� � � $<r��^��L)�?��� L���:4#�~MΈ���莆��]!��gs����Z�m4o�8��	Y#�뜥�xA9!�c"ܭn����m3QW��l2����g#p��\�,�n��B�F�T��ټ�hd��{�]حf�D]�'�j{4��K�����Q��,���@���B����cFe�}	�L̠�'��;�c�7�:�E��u�&]=R&���iE<���Gb��A8���0�u@&�-Ћ��sbΏ��>�]2��yqM�����R��8N�:�s�=��\���x��[�:�	}�~���Z���g[^����]݁.J�E1�x��u���N��pG�\�m�v�5)�ׇ�@]�	�mJC���	#:��R.����͐I��; d��5��ۨl��^��#�Z�:��5��p�SI����.게�Y�J���Z�\���gD��h�ez�u�(ap�ȶ�7A�^)�Z6,b��,3ZG\K&f��^�R)ӝR��lQUݕ<���;�`������Jz�48�e��5�S����*/��?R�d�zH����cJ���k��g���E"'&X:��8X_q���peK�����ֽ��Mp�S%�e�4�d�kO�M�n��t~��K[tO-�hS���2���Z��f֋�9Dʐ�&�
$�?�4#I�	<������P�>Q���\�E��E���f(t����b�W�[��\�M��Q����&(% �T���WbX?�K�j�H����^�C�'x-���d�.�F�C����$�L^��u������q�Cw����>{�c"�<����?�v5\Yu.]&RKTgW@��?�/�_<��*\��wP�:��YS�I�R����NX���������$n<��J���c'�b��P���#*S"1��R�8����0 ���Q�U΃]���Bcr�ɂ@\�d��K!��˄��/��/v�oo����d�KƉ�7%�UZ�Uz|��p`�pǾ��,>H�9�T��í�N�ֳ�l}������q4�vWg�� GF��ZѼ��Hи��)�l*t�	�2�T$�ٳd�D��0�#��H�O�<#���&d��r��x�-;��� W�U(gǸ^�H�Z�e����gxa�k����g�Ӽ�`p�r�v�3�#���C��Z�[ٵ\x�FX�*fVz�R/�����:�Z`/lw�|vmjF5dFgG^�L'��Rf0�����}��D�S�@�y��^������n&�q��l-��H���.���=��n��T�J(q-���^�ۿ���̂y�J+������|��=\�(�E�$=�tG�����m�ض�(X����L��&m�A�,�(SV~��15��ĞP'�ˑ��m����z�t���ݑAց��٬�Z��A9�>��fE�+�s �]M�L���w�a�ΕI�+57�r����ҡ3���4�������e.v��F�#"T?{�*t7���"F�҂AE�et}�b��w@�e�P��W����jzc@��^��S\T[���S2�&����b^N��#,��q&�
z��'82�:�al�����h��y�I^+#�UCΐ}Ժ��������Ԇ��D�P������X���T���C�&\�k �{�<��>ZL;�7���8�D���]�=��I=Q��nb��6	�+JI��8Co�d��~�D��1�y��U���:����]'~�x���1��9MN$@����R&S�&	�O����*����lxL-Vf%�<��-b�@�$���4l�KL��Pup��6w��b�$ʭ�7AL�5�ɾ#�p���ɣ8�ǕГL#A�$`_�����mo��8�͏� b�A�#��E����$%��!�x�:ALBB���A�cUk5�����u�*�ٗ�5BB�����0@ür�J�0 E!4E:��Xar�#by�Dt<��>h#��Φ�j_i(bν:V?�_�A���m9R�(�,��L���9��v�x�#&ܜ��Æp#,�Dޑ AL<�bb�.��:��q����V$�eh�zPIhy�|����c��tn����hD�P�\P�(%��W�m�r�Q�h�9��6��Mw��*�"Kς��9ps��lT�����$E����=��9g�]²K^rTĬȩ�3�z�;��z���g>����`A���K�]6��ߤ��~�==��7���Y3U]]]�����V���Z�	��4{�_T;N6W��=jFN��XJ�`��2Ɔ2�j������k���ڤ�-�Z#b�жI.�2�38ʘ��Y�V�~�|w<��H������d5&p̄'.N�ZBT>V�� C��ڋ"�h�-� &�����#T��lRK
$�~u��G��j*A��^�J�g��)k3�E�V����*��J\��$b�h���Y{�����{�,�X~q$�j5�-�ؐ@�d�<�Cj�
���|�.u��>��ֳ�(h�$� &�I� ��Q����1zV�|y\w��ӫV�%���5f4���#q쐮ex�]� b2�6i�7�C�`1>�ۀDhS��RT�hK����n�.���ɩ� ��FۢL���ߚ/Ƣ�'{�M%~|
��Z�<������������T����8�͠5���P��D]�Dn����ԉ8�i98�E����&?H�M a����紴�YA�?���3}���r��8�\�>>��� �Z��G�����h��m�	Q�M�w��-�5^�[�Ө����ܨ���<���!����&"��Lء&�@�놠>d����ѝhwg�5d��3k�x'U"�V��R�@���z㼕5վ��rRm�&���Bw��-�j��C���m��]HD]��lX�ɓ��|��%����
9�̿L���E�ɓ��5h9iL�D���<{`���_���]�VQ�!7%jA�.l�)������Ϸ��n^e�;s�Q� #6N��φ5��'�6�ŗ\�,*�ة��eфH[h��Kǫ���o�ޯ�X���:�f~,�!����n��1��<�MR�+�_��[ת��C�qzϪiK$Ң<��)?e_ΞP����p��r���Oq��~[��D�>�G��AąK������}M/Pߟ�v:RB����$A�*(���B�E�ָח�$T1q��d����ܮ�W��x=���3��ډcY��'t�5f�E�#	�8\(�Y}0�c`�w�i>�$���W���m��]�^F� ���ch�C쥷�#݈�e�;�qA�F��0���NE��}X�ZC�%�I� ��NRXJC-��m�A>��1�7_���_���-J�B�9�I�%�le9�Ŭ�*��	��g�t�	5h�ܸ��u,��ZI�N��D�r������߫��n�5�ՖY� �6aF���[��zALK�3�*�3Υ���m��!d���b�-Y^�X�׶\�-z�FK"D���j	��D�q�WT/[�4����]�v:f��*�{�7��'�+^ys�^�V�rs�ʋl&AL;��K����=&Jz)IF�G?�����8֍�Z^���NF���_����ř#��mB�4�aqD�(�f��QziI�ՀJ�������;�t�t�9�ò�~�y9N>�g��݅�*�^ާZƻ��Y��}�i/��EFN�����Oo8l�7���4�2qQx�Qi�8e�s��a��ut��=�2y˕�s����^����{3�5�J������y��6��q���7<5K�	;3hۡ�0i�d.�Y�u*���)�"�x-�)W)vJ*T6*q�	j�
s����I�nF����~��|��[����F��o3�.k�����&�b�;��u��2�i�j�a�RA���}�T�w�4���ry���y�f������U�[Ur}���D�+��Ga������]���EX�A�µ��c���qΧ'��a�7N���v{��*�7�qy�h>��$�L/Rb.g�Q��0�6h��+�H�Ł��H��݀���$T�����'�,�Ə6G�f��8�Gbsv��݂ۜ�;��R�~>�<�T�N9�:���U�ڑs%h�$��p�����a��� 7=�P�Ǯ$E��=F�
/5����b�jZ����*N
����	�#㘧��T>�����U"�%ܟ�����)��Q+ceTܜT/^�8�4��c�zP���mx�ډ�ր
�Qa/�����K�T�>"&��m�VڛM�9wkHN����R�2Z���-O.���R,J�S�&#%,eN�p�-Ϊ�8�Nސ@�$�Z��\u�C���1��I�ې��㨨|�$�qjR��oh^��� F�0����8w����Շ�Q��ڵ�.)��*l۠����=��;@��0�R�;t��.*i�$k�A��	#Yt��C� ���P���0O�0�������y`��u˰�eN����3=�K�J�Fk�
ʎJ�<��{mc�����A����^��|��1	#����F�
��ͪ�ܙ�6ò*��q�fa��8a�g�s!�VhL�5�`��|�u��^X�CfYy7��d�H�i'f�r�dDMo�8�A�W����m����-�6C/<=�w,���3F|\�cм�1l���-ܙ-W�M�ݔ,K�K�`�4+m��rn�&f���s���W�Q��FTj/YIm[��c�-�r�Vڽe����`/�\�K�/Gސ@#� � ��H�Ր�޲���a-�.v�����������s!��Qs�(g�]�u�UX�ځX4�A�5F�S�m�Êi�,e�'���V`IX�L���:�ű�T��&V����J�x��)�G��m�q�V��vm�\G���T2Ķ�*>`�7� �m/�c����.�< v|�%��c]���0p�m���&��pę7�Sq�8S��z+4΂}Տ��T��ܰ�_;n\�a��g*�Ͽ���v>����v��ㄧ����c�	;^ر��v~q�
�!�8�?o�r�=����[Y�*�����E��\�)�[9p�)�+3^"�����?fX�\�?M�X�J��V��K.��(�b�V	a���-���D5�bi.<��T��O�rGqJ7o�}^�폻_%v<ʦ:M��^� {7���7߸�'�8׶�1���ƾ+*��#����|��YD8�ޅ��8�қo�6bD$�jL�1ga=j��_���ʅ�ݛט4Э�*��(��FDCQN���wZ��re����������G'�k?U�/�<d/	b�PnX5-,.�xq���h@����E��ݛ.�8,?gğ/U4�� H����hAi��=D�K��Av���%΂����0U���	OaZai��?�r ��@��-�A3�9�����F}��A ���{T� Jt�	��}�򮤬����*���|��c�����d+	�����Ճ�|���gX~��Kސ@�#�e�ۣ7����̐@#��I5.2�* A����TZ��V8�\�mAv�/���Ty��!�I��xleTOX���J���b��!�6��+ �m~�Z��*ay����J��j	�H���e��u�m�'���r9DU���Sn�ZR�yWR�j_��z��TB�����:f���u�.�]�=L�������'.�/��oa=��8�DRNLW�G�����fCǛo%ǯ�X�|_8x�˨�[I~QqqzԢ���,�v�����%5�!h�ZXţ\>���R���4�a��rW��SR���,�f2�q�cMd�ʉ��2TR	�u�Y%"-�xq�ă�m���[�J��g�\�Z?�E5�~�<��]k�Q�gd"�1��SE�ơ���5��m��3�����^dޏF�Z�Ԋ%�*y)��ՊH���!J���&Mж��qD��8��qmf��B������Rn�j%�*���E�1N��'i@q&!�6I��Is���GUHʥ���&��@���PK��Z�������^�Cq�ck)P� ���\=�\�LT|9����n'���c��`�4h�L��GX�jz�⦯w�s� ���ݫ��߸��Պ��4������8��B�� �J]���	���������=�U���~�ƴ�$�ꐨJI���j'H(�2DD}P�ެj��ͨ5q= ������^Q�Ժ!�=�$�&ָ��$Ц�J{���%ꪝ�� ��M%�L��.��'�F�� �J��J&"�j!�6EDU
�Vʹ��jI&����JA�ޣJ�`�m��
K�)��0�K��~Tj��,�P��KCq!�6�G��T�0�붒�5� �j��0��r�E�3�t�R��z�*WrL� ��zű����?	5"h�Dc��Pm�p���Ҟ�8�c妐��޲8��!�G��|��\�bz5ܤ���/h� Ȧa�@��gA�8i7&��N;J� �jf���?�~q�ݟn"�J9��ǎF���)o��G�zO0_|��0�4�ROy];o��Ǜ**)g��`�����I�<ϳӻ�lH~{�M�kV�L�$҈ H��a� �*�q��*�L�r�Q'VO���=%)AuMI�
t�����v��
+����q\}��jU���ǫ���v���2&��۳m
+T<��r��'M��[޼L��Ǜ
*-g=�WUek�r�86�g縯�4�h[��6�ZDcBm��f"������b�[���c.�,��t�R	W�?J�&CAu��9�Yve��¡��U�F��(�4�ճ�ڏ��f/&C���0���ӊ��A�PL���/�����Rj��n�~� \d��VZ2l��a�'MO���ru+�{$�&���H�ZyQ*��g���#���h0y��
���U6|�����+�*I=��D#ԫ]��8s;�t�0bL�IBV6D\�ʻϴ)��7���W�2g���c1�n+���#�0���T�.�8�|N��tE�Yr�4/��c�J"x�ֱ�b2��1xj$>����ƺ>JC�H�i��x>��r��cn�j��o�0�$Ц�0!�c���2i�r�®�~�u�Y<�y�e���PaY�����څ�a)z;�/�tA�/\���r�+�b^�3F�i��/�#n�uX�bU)z�8i�/��-1�����OP�*�V&'����?���Ae��Vs�Q�5��'Pzq~���F�w-�V�L����b,m^�y��ʎH�VN��{F�˨t |T�J�Y�t%�*Z�|:-N2��3[U8�u�O<s�����Hd�����[�o�\L�������n��:�O7�ܔ�f �8mg��a�4A۽�������/CP8��F���IX���%�La�7N��r�9~ؽ����.���a�Ža�t���;Ǩ2���|f���`55���F~�2�]�����[��.�,�k�PR���r�VQ�H�$�&�J���Yi�YAU�$	$� ہ����-C����ϊ�Am����v�ϳ��%츼/�	�O���f;��䗱?Ӟ��t�ak�m���K�<U��}����+������k�?vPy�q����=ξq�G%�aX����)C9��e�c��	�vN���8Ϟ���J�!q)O��3����cNJ�ą�u8��d��u��/yK�Q=j���.���r�Axm\�)��x��B�\
������[�����x�#NR|i��P���*���0O|T3�Jtx_�|۽��,~(Ay{��u�(v�r��%��y�AqAa�r�)w��m�I-~��kPM�J�S��Ct:մ幎����@�؃%d�tD�c�,F���a���Txt��B���e�ŉCd��;.͎��ő H�Mq�{��_��.Ǚ���5XU���_��[������u�����է�kWB�˦��Z��_5�T�&.,��rǬ��(�[Vr�8��w�Z�&,f\�4�����-˘8�-T��Ⱥ�`a�1t�k��*�=m��=`vj�
g9%�,a����M,�|JS�r�j儘���BT�̹T
�n�;�qݵh�֧������ӭ^� �E��PA���	W�/́�H�|:�}�
7������ȭZ��jH1�4f��s�EZ�g	��hAAAu	�w�D�>��;^~���h�;3���ש��o�	�l�hvÙ��P֥��A�.xGK��-�ıF�k><�ܛy�y�
ټ\M8�uqtz��,^'��������uâ�3�������Ϫ�ĵ�?e��$��f�����P�쓙f-��\���!z�����0��''1�^�ҡo��Ey����7u(и;=�벢'9��nd�p�G���O!řiW�vf��?�~���
��X�a�W��8{�� ���`cz����ܟێ����
y�[qt�*5&M�Gs�\��\D��N�����v5*$�H>��>�`���#?�D5A�H��4�c��h`�����Ld�q��haO2h����=5|ޅ(��ru��u �59����)�:hs!e�3�C�5��ߍ^͌cN��",�Y��������^��ߋ��U� ���v@ADQ�x������W���z�G�C,_$jf�8��5���Fe/�8��zZ�-���`���^�w�+�[��AqP��m���J��y2�_�ZU��=�T5C����I�m�S�V�k1^���Qř�.��`�Y%�;R��;ch1��|��r#��_������8;2D�AT��W-�s��Z����q��k���oDk�Y�Ɇ#9ӣߞU3�~av��v���h���U��W�|�n�'�Vn�1� j��Mˌ����ؠ'���#��o��x9̂�	Wz81f��ɑ&�8J�Z�Q��K�Em41�g�߃���'���m}ר�����AL[��7z��̟qz�q���,�������c�q5��GԃV�)ǜ�Rh��U8�����<�gH�11�	��~X�櫠q��h���o�H/:$Ǥq�c�G���;<�[���u�a��0w}3o���d)dps����{̒��B��F)AO^H���?�Ƿ��zSݪ��.�jW�*~��Lc�K+�@b�^�^��m�2��ȃ b�~tB����s7������3�Fv�����=���:��Xx_޺h��;;jr�����s�]�z��j�Qq�<C� �I�BK�W�-����U����j�������N�z����?MN
����0�Q�YuT�&!b"���n��2��i��NdW�Rq<���+��)j�[�E#$u-��?�ĩP�݇�z�����-�a��s���c���$b�6x�xM�;�
��y"������+�T�*'q]��O�V�"�e2H��Q3�1���A�c�FD���H��6�����f��I>�V��#qxR�m�P������to|d�)�9�jfAL>��B����=���f`^zr�@3X���Ջf`����v�E�G�;z� A��c�89浳��Eb�s*jt��N�\��D�3�$6��̳�ۨh��c5kC��@#b�h��͖gq0ҳ��rf)3ƺh��M�J4�Þ$�[����m}D����718v��)�:�ܵCE�qm�
����APOAm�ZT5(��-1y+���>�Y�!�<	����I@������G\�
o�;~�ܔ�%�J�ʐm/�L�����c�iI�1�pK�p+��92jG�JN��\fD9H�M�\}eT\]�n�wkqww�����)�
����Stp�)��p���}���}�9�{'y����VPbj D�Gf*��G<�HͿ��U;�Á���(x��|�2��{��6o�L�������Hݝ�(ߩ����v4��T������^í�a�Œؓ�=���#	�W5����mgM���V?D�[+���^4�<��G����c̋��"�	�oZS�*��pb0�C��9����{����L���8wI� h4�Zuz��/h�VI\}�0��2��:(���ASiz�����0�	l Z�o�sK��?��\�%���q�j�D�:}���)�M��Pl��JJSO�|8�΍���[XŹZ7��m�x�>�T�1:�����rm ;���D�lY�Ć	i�1%_�U�p[Y�/���:%�H��]}���)�T�٧��\=�F.����P�p\(I�4G1ؓ�~n���A�T|w[�#��b�������,z/�rݓ��W g�{�%R���1�q�1]?�.PΞbqL�Y�gz�y���k�7�*��G����H&-w�0m>���S��(�
0Yl�JU�X}��&Ӂ�&�v�N*5���@�'F��d�a�:��1/Ԫ9�e�|z����~��߁�_U2�5j�Ui�%�ƈ%��~Mɚ�����u��k���ǭ��g��Ɗ��Ɏ���r�H�1ۛ�1�Q/�pHx:r dɶ�C�D�$ۡ���^���I۟��^W��{��H���3�rW8ne{��|Yw.���N���M�m�I2e��{��0��D5�s��R3�
�.�{-�b��c�;��>�Q�UO�Kտ�iA��2ţ�F�|�y���Jއɨ����^w'x�֞4s�:����K~�1���dE�ł}%Y��f]z�g[8������Q�/.*c�b�ж��Y�c�9깡�Fm�|��� �l�d��==�y�J�,���OW�!CL��|��;�F��w@3�sa�^l]U�\2��7�rN��x�,�øq�'�[�������ޮG��=�ŏ�?=)\�K�m��!��R�?�R�#��gJ
�V#-,�RN&};WbS�?H!�֖�o�.fY���Q����~+Z�j��i&S��г����>��70��@Aρ2��g��gS�A!�_~e���LYH�f��J;�{�W�@U"�L��AX����5�b��̗i������y
��[���Tį��j\��8�X�.j�3wՆ��k�9�:<��l�|8qM���\���r��#�;_�W�q{���xq%���em���c�cΉ���fm��,�sV�����/�=C+w:�1�fZuA�YV�w��N���Ew�	=�s��㪏��FA�A�-**�BLR,ZU^�2Y��S�e+S1I!��J�Q�vZ'��?��3����M)X�}u��]"�O^��m�l�f�f����&�g)SΎ����=��p5p��Q��ѻ����d��)DR���T]L��@�or�;�ۭ+�3t��8��v��P�%+��S^��%J��'�	��+�KD��?x��4.�^�U UQ©�3��rA��"�Sy�����(v�j��!2�DL5?p���+���۽3�#lˉU�aZ�LI��6<o#���˞����OF�����n��;�������yᲵ�ؔ����}6DV��\)1�,z�ِ[8V�T�,���d(���-k��U�6s�Ě�&��a-[����D勳�E��SH�+n_\q��.!Z\�i�}ۄN�[%�D���W��Hб���}I����g��rF���C�g�!W��M�+���ZU`ʚI)	M�4�v-�{��藌�EVv�U�j�����r�0p��'�( �R��a[��V\�bp���g�H�7#S�R�K)���G���:����@�iA���>���InO�V�c�����(������U���$���o�U52���t���5�%��)g�2?�)+1�%hT$YY�k^���6��{sm6�`w�nΉs�{ɟvX뢔����
�Dq�OQfY=jl�Ix�p�ꖦ@�E_��#l������Y���Z����K�UG
�۝3�ēW|�JN��Vx��d?�~�@�Q�uϠ�ۼ�S��p�䶯�\����Q�8�QNtM�AM�z��$�?�:�[h��ĩ�����4A��v>>�u#ːI`���v0�O,n��q��+��P�D�.�i�����⎵�x݈��9P3{���"�R>��s���#uͣɥ��L"���ҩ��~s׍���� #z�7��g��J����I�jH#�b��=��K'�����A��U���G$�"�P�i�����q�^����݇���aF'�<��׀
݂�?��29�� ��ek����¨��w���>Ͼ$���.F=�������A�QF�N�<;����נ���hmo���F8����[2�*���k��e��p��ͩW���R��(�`�����Ռ��Φ	,v��p��Ap�o)���_�׎:u�y:�[YچD��8�����CL��`y�մ�������؆Yv�]߹��~�*cK��<k�zѮ���S�^M���mꟍ
ЕJ�}�X��(ԀY~B
_���[|��zR�=�(�LO�%�Nr�P������؝4���Qv�*WbG�)F8Ę�!���o5?W+q��^�0�.Ւ�R4�m�Z�
��{F�6�*�zy�y�{?B�q,��s��X3x��@̀���ŗ�k�˱����!!J�c2��*��=��̛�p��Ù�*�fқ(��C�ɢ����bp��}��"{g�Qy@�Rդ�F��il;ȿ��V; ����$�S����!UB@Z�.���v��%e�s�Lgb���$�Ԙ�O`P����WH�����<�چ:��l���P��L�c'0�P���ѹ���BL7:#�/�����[��[4���㟂EP5����
��L��g�,RRQ"��S��f(���Ԩi�ra[�4q��ǅ�-@���G�q�m��<tQ�K��8���w
��\i�4ե5�i�Ks�5ш� 	��� �Fp�w�51��p���Z(��>�����vҕ_,�+����L�O�SK!��;޻�D5��N:O�`���:���.D�2ȼ
�ب�V2Jι���sM�'쯪���zw�x��Q6�idZ\&��/��Z�־�(P�3�=�al�tjo�*�io���������8����_�k�׃�	Oe�a��x��(��;�� ^���7|e|Ku��[���7㭗9N��u)�O��
����#r
�F_��ުTJ�䑰�&<�1�^�\M��$-���%	�㶜�h"2L�����=�K�/O�����JGm����n��}��[q�J!��A���)w7\�;Ltk߀<f=�g�[N&�W�N.�$����!��#�!*o>}F�^$�����dyWTY�$[�Gh��?LY���r�e&��3�-;�����#���%�)��S��b.�I+�EBDo����F�i�������l�<�$�'��T��ZU�<η����.����⅑r~ڪ�v1���� ��6S�FœC��=I�"���|���]��~B+mȈ��{�9�;��zawC����u|C�����S�A��ģh&c�x3��S�Ə���
H�#�(�a&���Ι�&~; � 5H�Y{KU��;3����&r��B�v�G6��6���V#[�!��W��-�T砖$�]��t�yH!��2�`r;�=sW�Vp0�L�B� ���DE+����F�E�:ú�"3�9��Z�����:�]�������P�W��ؠ#���U![�*KY�����t�����R�\=��8���n��%�y��I5��V���'�޸)�Љl4Z:��تG�q�v$���H�U�A�Q��n�""��
��Q8��g��F�B�0)�KP�wc�������O�[{���Rိ5�|�>ס@=���#��� 4Yk�|�z�$�+�S}ëN��m�9�K�.C�#ʠ�8(��jDN��샗U��]��ҡ:`��.s�m$m����V��n�r���[������B�}�$�e-�,�0\3"�d7D��Zv�ِ��Y4^t)�.�Mr_6�7#H������&lvl_�tE0�"@��(
�Ê���GI��I�������@��+�?����W.��VR�gG�c�=w�k���/>�-��t������ؐ��1�F��*oX���A�z��>����-��rw:!��V2��(�'�~�l%�dR�	}DV"dl�.���(�Y��O:C6O�%4�gtf�Eʜͱ���g��7���I�n�Z�9.vҜU3W�Q��D���4"6��ZP��7+����Y�L���N\:�<���)1��}����� ���*'�^O��2�1v��9p�nEzݨ�͇��ƅpXw��+Bϟ�L��Mv��?�Py��rŖ�*m����%&��w
��bJ���P�	�:�|�[6���6.�5����p�ﾁ�ڃOe q}�9��';/'�΋�h���;
��t�f	��>i�b|0>ô~=�����k��M7�6���y�L��*�pi�A�t4ƻ�q��۝a0d�=I���dP�&ו��/Z��)���.:-�ᾏ���h�cI!<}x8�*m��p�l�as��>��D1�^2�̔<X�Z=c���V
����
�|������{Ӏ�|v:_I�<�Y��>�?��(���	��V?�/ִԕBzfSH�.�7�,��kZOe���m��e�\�@��Nz������|����v��x�LÐ3)f��H�Ǡ��`��@�G�.�-*�v�;d�Ƕ�Ts�1Ƴ]���y����s|b��M�\�~�aW�'Bl��E��	���Y��V������͇-F����SnG�}�98v��ʲ�,�Z@%���Y�9�[�����ma~�-�����e�y_���-&>e�3��
C�V���u�[o�W(R����?J��V�b�x�tc����T�~��Y���j&�e�p��E=����<+���!s��s�Os�y��?��Uu��T �/a�[!���Ӻ�y��^7�w�h1)�D2��Nc]'�z���h�y_ E��jp�@y�:��@=v(g�gͺ`sbNV��?��.A`q�mg�ug�F <�:jOЉ�Or�o���d<[D8*�7�A�9)2g�ůr��S���A|��#�!9�d��FiF��d�*߶&�~����;]ǝx�S�m��x�N)����%T~!r'����swk{��,4��3��em�)RD�.��O ����w�����GĿ����ov�?�һ]�0�5��3)@3NP�E/
~$uZ_�8j+u�}�?���Z�d�@ߘz�gV�������z>H4ׯ�S�����I|P��Ƕ 뱬d�M��=�ט�����z՟�p��9,㖔Rl|�8�����@��_4��;�7�Κ�Xt�ԫRA�j���&�T(':^�,*��˃�G�"�;�7� q$��b�7�yL�q���B ���^�,sB��U��h� ��
l�<�A �w���z�LR�`����VV\�֔1f#��|]�����4k��}]�I�4�S���6pC7΅��H�g�:���Nǟ��f�N.��GU����{��@ �zN|��mFI-�U��-�C�n%�֮kh"�Q�:K��S�0�pV�D����M
q�������(�r��qׁTd�K��O� ����5府�
������6��C5�s�P:<�M��o6_Hc�$ �dD��#=��G6r�J��ʨb]t�46[��AI-2�eb�3�D��FH]���y�/q���K��Bk��g�L��v����8~bm��k�UUB�BIh%�<�����5V����F�D�Ol��9����<B��"u�Q�3)+�-u��Dčx,j@����Ԧ��X��eE��*E�~�z*#��)!r��8~�m!���p�D�z?��!�9�Y!�B&6����mY�� ٯ�a����U`��TA�
uoH��k+�n���[��g�,���-Z��<�8j2D����Ws*����f�X:���^���g�b����p�FT8�!V߭�6���h�kGʝ%�w9���y�Z9����	���;���MU�M6z��%QNX83x��oߛJ%�i�==���㖣��+���&�+K��v,��GJ�o1k�ǩ��e�fmV�%<H��`
:�>�J���w�{�rSq�oH`��5T��k�������2k��7K;E�X�d�+D��6KT5 ����^�n���H���ǈ�����>e%&�Ρ%"	i�YΣ[�F��S!�������V��|��ꢹZ�6}[13�*Cp�ik.�^�!�N"L�Ut����������F�O��ȑD�^|?�V��&H�{)]�PA�x�.E�B��l~���@�)�!}����a��6p��Z����)uCD��v�ǉ�Ɣ�l��_����5�E��>;S+Y�����k�*Mƌ��(n(��d�g��_�}��{�AJ�x�+s�ȷ_0���(��ֿ)��v'ב��I0�ʄ�î^TM�G�s�N9B��25�f}��U��� ��ml���~��)�,�6��_R⦿`���j�?TJ*+����ph�HD����C��&�4�Jg�,N,rKݲ�g��(Ļ��ΒE-��4$�\ר��Q�Bv~�Z��ʉ9�í�X��|҃$b�nzѰn�ݦ�Y�]����J����9���'��yN?U�`�����-����0�i�aQgsE�̧ha��%��, S����}�AO����XG]��C����!O���a �f�홨��or�
+�Gl���'���R�m��Nmf�z-,�M�ك��*�Kݹr���8��Y�ϋvJ'����گUVeYp����A�>hp��p��ZS�d�a�u��01�ݑo`��tU��ùxz<w�^�~�]G [���G��\U1�D'm���۔�!�s��f��U~����Iug����H~�_��xנ���%B%Pv�9c �a[���}]��_��:�t�~?`�K ���\������e^1 �X:g�r��ûuj��!�W���/b�<
�ݛ^�O��m({�!���.s̝���w�������^��QB_���kܔ��=;�G� Mýg��"O5g����8�w��	'�����[Ŏ��+����Qzm02�6	��J;:j����c%�������\�]%%�C#V�K��א(�1ULR���q�IX|���}�]������5b��2��,�%7Xlt�L�H)������9}G���pK���#�o?mxے���~�����W��X��W��"V�
�N;}�tC�:���k���K�3W�+�3h$J�=�蒦6�ސpě+f-bܽ��dɭ�y-��_��>�T�O#���|����8��y�.���;�N���<�jB\�9 ����\9���v��P~��Jm�cBf ���ay����[�Dr��d��X*��ߥ���^vf��>�2��k���.qZ���H�mW�渆^�DC�g��+�Z�g3�֬!ۍ�"�͘�Gwn�w~*��#�;��̳���Խ�u1(tĢ�O�Bw��P���z�p��-.�o ݸ6M�^��@���/�^�;)I�v��BJTw������kl�G�w���w��k�j���җC��ٶ}��z3n�b�[i�LuAt�V͘1
��6��&ۇ�O���t(�,��c�������?�`R��X��,T�	5�a�}'��(��e�_N��&���;��O��C�_/#DV��^�����"$|'2޽�ī�[74א��zMN�z�7������mң����Yv��T0d��UI��N��
ƹ���U0ֳmĜ՛���� _����Y�H?���>0F޾:��j�G�ȁ����>�*^��)L3ᤑ�Y�9�K��l�؅䱲o�#�ޔw���3�L����:)߉z�������٫�U��O�y>��s^Q�UJ��5���/�qh͑�=���5��K'V-�v<wV(�z�)ur��sc�u��\�[ݝwGy���5c�����#��0}�Dg�X�TT>��`���b���.�����3��xQ�
��J[{r֓VS�a�zUS�)��N�ƻiV��D�����ͧv���N���ծ+������޸�Y�y%�]	�zDV<K�CQD��`���{)"��G�r~�����4�� �^��e�r8t�������٬���ܡ�Z����x� ��C�X�r4y����2����_�h.���7
���I�O\�*�7����O���2c �/��s��X/��6�j�o&)?�'�E�����X�3��rq���P��5��gsNِ��鱶�S�9���!Q�
�8F���.ЀuJ��"RZ��P�/���n�-�����
=���t��I�S~��<�b&�T6?��f6i�z��,*�F�����NX<��������ͤ7}l�n).�ާ��Jm�y�fn�i���ӌ�@�F��0Ɖb)t/z	��w�ysپX�)�v����X�Q2E;���$ˢgt{~���z��'Z|��N+8�!
����Է���L`�[|%��|CCI����m��;�n9��HV+u�BD��!�-ht�AC׭�i��Eq�H��N���0P������L���v�j�(�8�3�����c���� (�ƔjQ���fO���<�A��T������m�|
����oiw2�M�NrQP�e��R�U�B�u%{I6 cfgU��4_�����چsh4ɼ:~+���p.G;��L�f���(�¬���J�hHN�(ehzv�no����E��T�?"��l=�2d��.U$�X��P��HkkA�h/jMjZ�Dۀic�Z�x��`e�&=��Ӗ���u�e{%���9���%�M,g1�9BĔƜkp�y�g%���C62S��
�h@����P�F���M�`尙�]�qF��;�S?���/(���>>���f$:��$�o����_j�Ӧ��!|Fym����{9�g<�e��6�PK�^��L]7���5V`jͱ��߿C����xv[9�jU�=#��Y߼蘳s4i�϶�F�l�ϟZ<�I����Ź�d��%�M��,�`-.zqƋ�d�rZ�m��lr���г��JT{�p����њO�k�>����wJ��<�*�_{�x-G+w_q^���Vg{©n�_6�DL_����pVO�U|�wX> 9DQ}��eX�W�"��{&P��I�]ԃq �C�hp�%,:���3�?�����J��|�l���:~�x�Zg���!Y�z�{V
lL9�3?��3�K�D}y��b��������F�"��x�CU����na>I`g���`�gnE���gy�b�_LOB�����*J�Y�����L;{lJ��g��e�r�ɝq�X-��w��lCY��޹.:���,5�_OJ������6��Qh����\C}�R��/�n��;	�r�|���Ez�y�U��Rδ����2��su��0ɂ�}��q�W�ļ��`�kf�g[/k�_���À�9.�Q��������}-
|B[ 鵁��9υzͮB4f]�x�Ң+�y�vV����`������ws���5�.PxR6� ~k�e@���?��m��VF��m����!Y���������)�a��9���e�ҡ��~Y�ah��6�#�{C��E6z�:����8�vߓ��{���gk鮨	�l]�uI�
��>~&�yIu;�%X��!o��h���m5/񬾅pi�Z��9|^�D)�h�:��l=߰��E��;e�����廩�/��F��y�n�,m�z�/�����Ŏ�0[܎>Mvj�r͗$�=oy���{��`�r���"c9/�e���ؤǳu��C�/ �^5�Qq�>����v�{��ESlg�ǚ9c�8,�%T�SkRh������w'�Dq�J����g�<i�*�;O:m:�h{ͪ�}�^��9����ҏ�����k���F�����f5]��mj�i��k���ʛ�C ŐU��%}�+[��	�O��Y1^�~	��N��oe��'镞@�yy��͂W^\~um'��ͫ�ӏ{���y}��u�L�q�{@�ʞ�Q����Q�Nr�7�q��Em�P�3��F�C/��x�ıigH�nG���IL�7;F��҄�BܵC�w�����(ڠ7��_j"N�r�����r�K��aV;=aM$|�FKU�Ȕi�i���c�*Wr�g-,';����ȽM��U<»)^M',�BM��W)I6�G=Zر(H�y�����~>��r�~�虬�-�N0��0�RV�jgΡBW��Rh
D�d�قw�hE�K*Ϯ�o��$���L�j6����yq�L|]����x����H��^,��D��q�k�KcKD@!LH�Qg��A�]�n{e�i p������ ��~-ʲdt�{M"F޴��'6�I����E�<�_��b�LwKc�s�p�����_>e1��/�>/����'*�����_abm�6,'��r1��5�ig?���.� B���$�D�4�.�V�U��,�Ǧ�l�)v�-��u�b�DY�.ۓ�1W�h�C�>{G9���8��5�h Y���PV���<
On\+��v��j�G?SƆ��Z�5oW>���xSw�����UC�!�g��"@y��D��{��UU��@��u���mbv�st�]�?_�w���V���{����i�H���q������_�h	�z���`�H���@~�ӱV|�*G����L�I3���Xw�7u�dk������
M:��%�ա�1�,����8�
�9�t�`~$}��Z�a���0��H����_�1\|�	�D)�iP��&s6�������6�X���!�		��������Ͳ�p��}4����Ƴ*bG�t=衏�~E��2��������[bH[ﰤ�#�s�	&���ñW��5k��q6��ϯ��d���~)���Is���l�P�����l�������L{y,�XR;�7s����fÉ��e7JtN.9���6G��b�$�ޛ�h�w`�����S���˚���}�K���M�R�z����<�T�9����4�E=����m=o)��:��ZQ.T�Ҙ����X�H[�?�u�jؖ�	+��Ć-\����ɋp�5� �0�_�YT�`�����zb�z6�Nb�ي������!j��t���}L,���Q�\)ږ�����RR����콻�g�z�J!ʘ��y��4F�w2X !OK�|?|��C����í�n{�^N���Vӱ�1S0���K��ʌ!��a� �F���5+)�}��q8�(�if�p-1����$ӭ�`��	������⸁����3ՖYՊ6R���"�5%xz�Le�ۆk�������RP���F��,�,�sԮI,�b�k�d������+3�uax��<����4�C@%�*M��w�V}��m^�U�
�~B�e�{SQ����N ܒ���w�wrD35�3��5�NӤ=�8���6!"���*��zҗ��1|��[��/�oe��	\"J�@�PfC���}�e�V�//���?�9�d>"�}�������Q��m�ېd�!nDѯV5��!*����F��&.�uT�g�?ٗ��&Ԁ�=����c�1D��[�K�j�% b�"��:X�H/�֬�pp�1È'��<���ȪX1����҈عgh��osf�(��ahJ��:q�c��z�P���2&RS.�O$*��B�zYq\g����i�|Jb�J<31�^����S�$�W�G�-n{|&)g�s5'��&���l�[�)��)D�҇%��c�4�WCMd�HkG�#jG�<��؎,ꅁa�ֿ˚��xq���A�I6�۹�!S�tdV�݄v���e��7�Ѭ?h�9�m2��f}���G.(gtУ�ؘ�ʋ�PNF}�I�]�cN����L����˸ �8���FX 8z�UHx+��;&�*Sz�Ѵ�?\�J}4597)#�E:Nx��E�'�h�)F�V����/�!3�S<f��+��΄�J��%5�ƭ�����Ȩ�Q��7�T�zE�V�d��+��zoN��'��Ұ݅H�%�K���K�0�6���{���}�j��˵�v��Z��U�^�5\dZ/��p�i{*6�ӣک4�Tj5���������Xz��z��fNA&�0;�k��W�F��{Pw��)��sk�Q������T��83��9���� %���������ݶ&�(���13�y;�3$u�6�nR�4-
�=M�L>�%�����7���a�����s�QX:�
�#���-�!��-��K���yb(G"�ʹcZ�N�	���X�gD�c�E��f"��-
������0%wqe0mi�HZ�}��6�(X턔�ϡ7WόĪ���/�X)�i�Ŀ����ڲ, ݈#��9O��t����s'�s���u�D��f@Rxuc�L�<���֥m�<'J�(������%X�������������~��O��������+�ћnF�s�c1#�XS/�\��K�s���TZ���~�Tsa	��tr�﷖�dR{a7��n����D{��B����R-��W�F�b��?mb����hv0�'R�|c�=�xȡ�=a�0T�5\f��
f�L��pS ���� ��ڶ�lW	���4��U'���>ctn�L'�)#t�M�7Ȃɏr:����N�$`���/kw~�o�2���b?����%�&�xg����8��9��4ӌaQ]c[�������U�����>m���M�&��>ᅢ�K�"������@l6.VnӚ�'�ڨ>���vQ�����˸�n��T�=�4�ԅ_�x�3��{�m1cE?�j��F"�������4�u܏�������({�;��	��AKS8�w΁�����}k��+�0�$�_{��_p�;,�@�s�, �ҿJ��NFʓ�~����~��n���zN�[�QBO��{|�(��Ad��MTw����.��0�E�O"V��Omb5aMƣ �c<�T?�d2���~a�=��3lpp���WT��x�VQ�r �}M	�'0�����9�M�D�:J��
#T��6�1�oE\r���]��}a<��ém���)
`��3���"%�侄� t0�5"�m�
�%�в����$��jƲ�Mnn�uc@�e<�ԊY�>n����.��5Φ3��m���ԉ�<mՎh_�>�6���oڅF��Ii�"Y �D��?o�� TEǶ��a��r��������9s_,U�h��U���6Ӷ�E�NG8�_|P$e5x8T�P��E��Yq���I�b���f7��D�/��3T�-�'�V
�m���)q�ڽ�䩶U=̫k\,0�R���7��E
�'�y��'����ԋJ.�b��[.�ԝ�&[�V�<�\B[�:�t��>j���r����0��؛�?6�(m���S\>��g��o���K�>��V���x�"[u�Sɐ���˔�x�9��U���z���sK��K��b&`%PQ4�����3/0J;JLh0͆�\��Q�{��*��ˏ',�}_M���	��)��N�?��]w�뚫.���p`�a)٦�>X�{�՚w����_X����ì�!0BT�!N��,��c7��	�VG-�
��P�Ik�(T�aSH��1�B�*��X�5Z\��)��~�E��\�U�͐r��Ã2���8�P=�W�
I褎\�ڭì�`�jΆ
�Ʋ�~VD!�'8;�w髌�ͯ�:D7�2,?PE)����)1.�j2C��i�1��Q1�`߹�˷���O��=���5�e�B�D!�F�["U,�w@��8m��_���6~-7�H~�GTQƦ��ap#�f�N4h蛝�{a�rB)V�@�W<KX�6���W�z���rST�7ܲ�v�����a,9�fE�\��I�����%kK&E*�7�p�`�#�Q'�զ�i\i
kk惨�9�zI�e����+*tUk��	s�C�`�/ڹ�@S�k$4@��n�%]W��*���Ѭ�v<V��)S/�v^�Ư��BX��F�ԑ.�X�W��ģb���|7Ӎ[���Ρ� R�(؝�k̗�"6b0����5����v ��i�Q��b�-�y��.��hXȶsӿ)�<�P���Α��c(��4���H�67a�rg����M��RՖ�.c���$i/�m��Ľ&��,,�w�t�1�>��_LHM|�#�� �vd���K����0�,Ɵ���.��p�k�wo[�+�H
Br���\'�tP0��*������ƀg�s�'�"k�5���8:#wB�"��*7:B�pRr�[�DZNp�I9�$���8�yw(cT��;��w�O�Q�����J�D�P�����d������+z���4��KD�6,Z��h�����aDNgK���^�m�]Ni��a�a��v�o�q
�`�;FbS#S�g���`��o�������#�N ŉ?��3�z��*�Az��Q�^k��Q�5�c�������W����Ҍ�F��Gk�	�7o�G_��1���1E+8���:.�8��qs�k�$ǔp�� G���؅�\�b��#S6i��})@r������N�}C��NkI��ʷ��H���F�<�<��W��Fl��vq�X2Vp���Jx��F�K�hd`�����gu��0���r]���B]�ꦆ9SV}&�tiȵ�8���}%�-��i�+�/J�}5	g%���D˝�'+_/����t�70,?q��� s���),WK�Y9���㬫��K����"���G������b������?Pܬ+���%ns��K�DbT�}��_��}��)�����):�4}B�r=�W�t��a�WJ���X/5��q��'���C	b����:�g}9bRjb��fI�_���6���P�FlM�>F&�������Ȅnz���Q>�]��x2�s�R�
����L"'̑w�ҐHT���XR��`ߵ�.����9��z~e�C���N;1�E1����՗gl8�Wz�O��J�|9���oqv'��N:-�U�)�j�Mn#L�O��.+g��И7����}��$���8l�����9� ��R� �Z෦S�ܯΘ�\�f���Z�R^@����ap$,R��r�~+ý�Ll��UYNL����1r����:W���;>��fY6�Fqg�rge�<���J��_�?�ǅ@I�dGA�d.�kd�JF�/�M��[	O���,��tФa��:1E�����D�,����S9\��B�-�ӭ��2�s���t55w���}�n�t|s���H^Hʻ�9����
S���Ih��Й��	7��^v[@���W�e��7�_S�_=�Z`|�6���.�y�����&:��OTA�%��>c�h�,,��HL�K�}F}zg�Y4e�bσ�Jy���i��톑�
1�����}��B^a�����XL������-����Ak��2�g�ɗj��ȩ7d����a6���0Hiǻny��|��|��Y����zԉ����.� $�V��w�3Oa�����d�f:\V�)j�m�_k�;͜������^X~� e���U��؀Ε1�v+5v��6b�ͧ�f_W��6u<K���������_����8V7�Чvi-�{���T�t��C[��:U�#�;�VƎE@j�)ᱥ����\�8����V~�N��W[�Z0E�I�T����JclOx�����3���	�T�im67�p����ѴM����@�.���cp��+�L���ο<iG��%|Gj��o���D|�F��{+��w$�+`h���X��P��׷���>���R��/f�ӿ�Gc�r���ό��CiC����ُ������}��?T����q�b���Z�q�S0V��>J�����L�%X�ӷ]�����~��?[iE�@���V�h+|�vX������Ckv�
7ގ�����A����sf:c���1�Q܆����'�Iѻ+���~/�W��xjhv����^��P=�u�%������Q]��1"�����qg�tm�?�Z-� ۣ˹�};�� �`Ο�̶�0d����Ը��u���D2�v-�H'��Z�y�;+��q�-L]_�� (~�ɖ�1|W�jupd6��r�f�}�S�&�6,�|0ݍ�ǁNm[�^ݽlX:�T�M>z�x��G^06n��<��,o��C���.����ߐ��)_G�m�����w�!�>�� h�\BpMp��\���ν�<݇��ݻ���v�Z�zW��4(�&q�VU]p���]��+|�Z��ֈ3��o8�Xu�#_9<�&l��ڽ�H��͜%(�'����Y������4M�&�1��]��܇�:�������9z+m��^n�O��D���/��Ktss���[A�I��_D#%z�R�$!g��������	~R����c��{��z~_9�%8е���o#F�=d�����CGF'����0!n�>sOR{��,�,��^]+����@�����'E����S٩��eʼ���j�c���8����Km��=B����I�g�������n����[�^�:2�H���\���1�︖�C�˽�����w���B$�bw�����+9����!�0�.B����Ϳz��5�b&��*��uf���o,��љ~%��Pc���Ϯ��)��������k���`ok��IvUhY`�K������St-��z�~�G�%�l�2�5%��I�p�EY��.S�ƉN�ko_�!��ǌ�}��ߗ��a
������d�cW�:c��V*��K���}O��G`��h�c�������!i��Pf,x���ו��dzZ�T���J�,bv��|^]xC�Ǣ�:ƺ���5DRǘI���TA��wХ���]��g���}�!k�Y�m��L��{jP��R�}},-UF)He$R��ǑټSHΖ�E�������I9��֘D�&�'m��\�����l�2)��������KS��`�������Hc�X* *���A�
�#�/��y-��O��w�V��K#D�@T��"Ήd��q��2ؚl¡$9H�އ�~&D,z��Kj?QV����G�,c���`�ӣ�$-�l�����=�#S_�^����ħ�O�g�=Ҁ�x�+0.����ҡ��R�n� �}f��HAI�����lї�qj�H�	��H61w�:���e�Q�+7Y�D]r��#Wߺ.Y�y��yX0#�̈"Ʊ$>� ��TH菥�o��9���q���˛r�,q�qqLIT�	���k���Fᩓ13\\�/�C	cA�vN=%��e�7q�x\��m#���:���0x�6���լДF��zP·�ȔH���F@;�&�SK|�ͯ�o(�rl���Zb���C�������.IG�t���%�T�w��r�ѻ�����Do���d�����C���{HS#S�l%��V7i �;V��)�(��wZ��&�j�%a�$-^8��./58��_��TShF���Y���t����.)w+&���A�Yd�͋�x{>B�k�:/����IŃ��؛1�F�X�b�U�/�DF�~����h�͗��(�
<t�a+yB��3޻֯��$B�q�������!�����1����L��hS��R�&�˝�n���lf�2be����K�CI�CzX#��]!��@���P`h���P����41&�S���y2���p�d;�}F�������KJVH�*'�h���h�m�N*����_��?P0�A�>_�g���
g�(�zv�;�����֬$�^�;���~���H��X�O"��}�	��¦vX�5��Z�@�< �0<��4)������+4!u��` `A!*��le���~H�÷���v$��|~���ǘ;U���?�\.eww�K`E֤ᑈ��l�[�Љ�%Kut/��ݶ�Hǲ�"�^(��}�2X� 'ЦÎ��}��zτ.G������7�Y�9bE
?z?V�d63&��7��}�
"T@$�c�0�8�5��qa�Wxo�)�Fj��͝���<U�ə��WX
��f��KŢ�7�S�J]S!hL)W̰�TWU1;v����P��omm5���5�)�wF3mX�.cq
"S�먲����*z��NL�Www�/�jj�9����d\S��' ����T ���;�#�������,]#����p%����� �mJh�("��@/Ճ3�er[���Š�vTM�I��ř�Т$�L�S�Ңw-�#e���Sm�����Y�^���z]�W�|�ߴ�T��a>�Q6����@�{�-(�ކ�c�� ���7��}����I�B*��f��r>� 5����|u]3jq���xtr�a�A��<����tБ���!�%���0v��g���@�o�P��%趞���6����;�9kZ��4-ز!�	�=73ænjjZ:ᤩ_g֭bC��Nk=��W9�4J������%ϸ ^�1��k�M�A|Kl�?�`t���oU�����̠_|�D(1rgG�O��t;��w\��_,fC��2u���UZ��ޥm<R�.G���g�J:ǝ�~!ݣ�P~�BQ3/�=kv���<_�sz�ǍջG[��a��1�؟z��l���_�a���E�p���m�!U���:!�r4���,���ns�ܒ�v�/�ָJ�������d�p�dA76o���8�!�j�
+�M��}k6n��nR��0��̟�U��hIh��>�U8d���k�Eg�mxI���'�7�ۭ�����jI���4�(C��r�{n����z����8����"��i�sԉ3�������NRV�.�u�#I������� R�d^ρ��q��Q�0s�Q#��=Q���.������ʆ�Ԅ�1�#���� L�|�a}��N�ʀKr`��1�C{�G��-P�Y�l�Z�h7pX��Lyv��M/�����RD��4�rn-L���jj���k�cf�/Âa����7%��KA:��|r�SC���⤌��|���o��t��\.N{l������?�(_�r���x�d�?_%G�7�\y��:5z�J����Uc��j'	Mr�������H��� DB����ϲר�u�q���I�Jŕ��n�Y�.�d�1��Y@�������zSq.�wϖ��t~������%�42�(U]��������]uR��f3�kz�q�Ka����n2||T�8�1�'h�o�!<ښ��⨾W��m-�5�`��F��Y
KK�:�L&��>	R;��綞gBR랇#��Y�����F8:�|���-X�����|���v�wh|ָ�H�E�fE��>��*�cR ���u(��n4�|4쥠��Qbf��Aj��R�z��7��-���JZ_ݚ��n������K!X��4n���?師o"����#vݠH�r�)�}@�U�QBFhD{i&��jm�'����P^1v�{X�ŉ�d�,�!�f���`(��q�&�Q ��%V�a��S�T�ij�$���}c2�-]dJ<7�h^O�2d��ZC��$*��!�W�5b"��`ww�p���n�N�vXA�z����s8�ju������B�Ƅ�u���������W-G�!f$�Ʉ�������Q�.O19
���c&Ҭ��]�L�j�ٓ����~�����h���ƙ����}@�^YT�C���}ޮ��R�R�H]�}k��������O��Ǟ��p����b��ղ�|%a�}bt>z�/!Q�f�m��&� Z����[[n^���r���;ǈ
��ka�X+��zB�LT��މ]r��U
�+X���\�Da�sh�ǫY5�sb�@%>kf'�΀j�lGڅ��J�Ρx"��o��S^$	9�v�����@��,U$Y�2�0"�G����#Rw3����M�,�ZD���|fB�u{��e�7JLmC��QY��EA:{�QP�ܼ���ہ��OC�C�M�H�*��X漈���[zH)��!aOϱ~�%3��ue�wfpjA�drkظk��_�p`s�|���^�7��hl����NCI'3��?92�a�i)B�R5o�mKOlC��B��ݢ�W�R��G0D����9~�!]�߉��$ИX�[�
�(�~ڍi6i�=x�Űd��ԩ�Q�ꁹ~�&�nJ
bmڲ 4>c_Դ�g�w$�Rp.aL��Kj�SJaX����B.e��	7���g�buS�����0D�ٻ8��[p�(���}>z�K�6��/!��QPh����*��=�y��@q��1KM��L���������2å�ìr�?��mN�B en�M���/�'3j�x�x����s'dK|�<�'�����O2h|�a�ȹ�y������_2��`(��&oQ��L�CMMQy��P��o��*4m�NV/��x�`3q���FB�~e��۪��b��)�^n� OonݖUF6$Z��f�[Z���C������2,�7cy�^�O��.��@VZ�J��WU�-T%6�{}�������6��~w�;>��Ћ�B>d�P���Sc�K�e(����nL�^ڂCo��j����f���|Hb(��%ەr��h�s���I7��)N�1����P-����Ụf
e��Ǐ`���'@������~�'�w��ҏ������6JB��ߵo��D�:�|�Bzl�*��P�y1e���e�;g��M��C����o�2-�����xjp2���^1wK$<5"�]�4��J�s�o	Q[�$QB̉?#k�	�)`k�9�qVz�Q�N��n�i\Z:|�ϙp�r!�qa5To�Wm�G��,���tD��$�;,m%90!��Td���#�>����|dc08g.����<@Xxςpސ�]ggg��������Hpnb5�PܫY�[�,�plog�ݮ�Q��<�3������%T����ĕ���d���޸����Eɾ$�dtx��̷�$m���{&�l$������`h���b4�Q����N6�Ι��;^b~qq���?6v8Բt�jjՌ���>b-���>�˯t��13srpp�L�F���q~ �ĩ-cjC!��8�Z�l` �WNm���x.���ʌ��s���v{�5�v�a�
N����J%�����'u����]bC99�=dL��<�\��b&�S��|au<S�e)�Z-I�6c�����-����Rc�ع���Z�n��c�/"R~���9���r��g����Jл���ݫVW�w?�+������w����9f]��;5j{��rԦ!�>�M4>�:�>;�-( o�����ᘗ���,���7{��ť��!O���S��O��~����LLN$�'����&�drY�����6�������G���M�Sg�:m���Q������ہ����Q�<3H��D�E�'oNVf�C�T�I��U�]����|�Ӕ|41��$��*����K?�R����ij�����8L~}xx� ����AԆ�`|5j5�����N����VX�d2Q�C�B�XHT1��S�?1�l��,���ռR3�g��K���iU��n�0��;�5�e����ҹ�9�F�������S��J��ɉ����-�%�B䥘����Z\�c�� H+��zڐݗ͏ �"ܛ���{%ŝa�p$�t�Sa�b�f��o{�K�3Q�8s���A��B���̇�<�YީSm�IsP+kV}<���L��0H���EC���Fl���A��?���;Y�5��۪1�:���t{�z���X{"�[�!i�$3�cۮ�����<�T7$<nn�G�P��{�j�+��#'�c�3K{MS��5��\������3[��r�B.��)��m�x�(�I�W���j���E�D�V2�]~�--mU@ZB ���;r�Q�#������|A�B�v��i�#���|sR'�ye:�{*/����������G�g��]}V"J.��PƵ�t���uE�:���{�8��ǳ���v��� n}lr8�0�+&�e��ԡ$7p{�\z/^�]�Nb��]M�ِ�|���Ѧ9�$�z�_gRxﲸ�ix�<�|"p��qpO��X��}�R��{p7��bG�lm���y����th�����\���X���%`��GK3��[8��A��@��e�j�d�D8C�|�x}d�%٫�����T�Xn	�T��+�!#.�v]�f���⧻-=�F̈�b7 <���x���'g�=��]��"L#�r����n#���\���D��K�Ļ3L!\g���^�$�(����p����.�'=�ڋ����3�3��gb�u�,;f�Kص����+���Z�7�&X���q�����*��h�����ݤ���D7J ns&�sKЇ��(R���P��S�RV�OӁ�V^��`��m��1�^!�IU������Y�f���6�;}7�>g)�_��1����t�䅧��c���,������ꄥ~�z���Y֛v*,��.���]��H����\����t�D����w�`�W\��@#NQ�	I�b����8�����`�ioȯ���.��pꈈ�`us���kU�g�s .�wH�Ӵ�pT�����|}s]YRb�𷆏�qsk3�,��崗�ZS��Ѣ'�3��n,Xe������"1��Om���$���DZf���3�����Jo.o��}M%�J�m5F���[1_{��\r@�������5:ͩ�u�[��J��
C`t�F�����Ψ���p�����N��^`/�+��L�(9<ۢ��)*/�"��|�|h\>����{�h�m�#ݚiRm���h~8�nzy�a����@�ͦg�mK�]|���D]x�f���uRJ?9�Z���l8���]�3F IWmb!�m�����bú��Q5<��.��[��q?�����J�U�败���������A��`��%�`U�[/,�"��B���L���-h��mj����e���7�?1��5��r�A��b���X��q��vcF@B[�'��T[~�lnYHy�Y;Ôk/-%в)&�z6���g��Z=!q1𫺦sl���3�PqڂI���u�޶�p[ޗ�C_v���L���U��aXE��c|�a�!��N�-,h���^*���6)��01���H���&'�v����7ǫD�Ņxv��06%qg�>/e���_0���+�σ�����g�@]�:��|g_�%�� �/�������v�%0�	1�D}���1!'M�/��㵓f�o\b/������?u�6��
=��ޜ�.\�H�����8��7��Uw����N�!�:�\�V������1;U�IN��{�T�����5�=q]?HM�K\f�n�<�o}� Do�y���������Te|m�G����L.|����zQ�qYie�Y�#N�O?�m8�2)�
,���=̿�o^��fk_��4;����a훻�u����m�	����-ܩ� *�VW��׵r��LEnfi���������S���!��-�w�_'�SG�Q���a�l��ń��ƛ�[őn�4V��{�r�eQm8��-�e�z����}��3���0���ɧx�|1����ukZ�Z���b�>�XypmI�vO���H:��XxQG�u���V���e.oWC��8��1��P���Mź7K�RKZ�+�f��P7��J�`��4�?�&f- յz��"B7����
pZ
+D������^
���l����|m��̵�5��@߳������\����C���^?p�h���T9����%��I{&�`������u��o���ʖr2��͒��I��wX�hY��B�Z�9~�'�'a�OM�Pg�]�
Pj��� $���կ��i��֎�^��\ƪ��䗁�>{7����Ә���r�o�B��}N������z�mE�
����!|��Z!�d>��ՙ�������2��3s|���'�2�w�gL^ƛ��@�3�����̀���s�d�4�p�8+K���ކ�[��<{}0^��tb�Jd�k�W����/O�%
h��A��}�}�#��%��~Ke"������	�L��s���D�b|̎�`�Z$y7T���9�|>9[�O��PJ��5FM��~~��7[�����+��Ԣ�WT�E��O^x+A�j#��z�p�MW[Q�(Q$�+�ɽ�������6tbi��[�*w��,t_8���[��:�֚8���Bk���� �8tX�7�u[��'���8��y�2e�=�M���n��p]��QU\窷��P�Xr�0�A�7&ӛ��￺܄o�w���z�K2�kp���Hib8{���LVn_nJ��=�-5���T��� :'��s���ԨC ���}A~�������K^n�ƍs�+���)"`r؞,:�¹_��b>�2Qn��C����U���A�U���z�5�<�X�UU��ʫD���K/�/�E�Υ�M�T���j(NT�7xe�;��&�dc����;Y�;�OM/$_]궏�qY*չ��b~���N�Mtf[��&݌��ְ�Z"���{�,������r��"�&3�xο��6&�
�!@���W;������fK�BH�m���i-o��j��:�jF��>�>�������;P"g�̎���$q���'�t���w+{�]�d�77�<o�Y�˹j$&���2y|v�j������EnǕ���\KdT)f'�ќs@�T�������?��b�K���<�.@��ͮ+���b-��yIi�l��G��Hhw�"/, ����9)�4Nֻu�-��o�T�JSy�7��XR[[���2	YU���-ᱚ�%q��1��7F[�U1��O�93g��Υ{�R�@{�J�������zue��$a��bS��y+x�8LaX̽b�B"��y���r%��]��}er�^t�<A�����`����&KN�a��vC��
���bnrA]Nˮ'k�u,�����TĥD�6���ⷯ�(�9V�J�&�
�Xko���F����VZ]�{��D�B�7Sd獫��	3p�����3��y�+H��M�Q c�)ʡcp��m؁P�M�B]�͛p!�S�9PAr�9������ۑ�fːdy�US�9i������^y�pv��//sLhk
{���_�t���^��Ř�Ѥ���2�3l�{~|9�%oy��a+�14 ��2ւp�:&��9w5n3��a�.��a>���V9zN�\*5����\�{Rm{�<Yq�J�~��U�+Ӏ�	�M�����Q��.ԗr��WSS�ʋ��/���؉���9��'	u�D�}{��Q��c��l�w�h([G)��K0T	�3X��cː����� S㇇SޗR���`Ep��޸+��Β�I�� ӎ��pjf�{���yI0�%VAA<. ���;������{��_���
h`rM	�1a�4*z�ҰB:�=�)u��+��z�eug�,�����JRE+!0P�AHz�3[���pxt�3�V����q�~4wW�h�Sz���IFB�m|�ؼ�)�=4��Ps�r����Ebb\�DT�E]�Q�v�l�V�=�R#8��@�t&�E*X����~g3�d@v��lJu�XV0��Ћ�NfY�Bh�ߞu�Oԫ����<�A[���R�C*X�X1Gp1V��R1���mg�*�iIh�\��>ftL�G:".����)t����_���5<1��!1n��K"����;]��+h,z��e̛#|+*�p�]���������1p+q5)Y��2ߺGB�w�i�s�n�Ro!�һ�������m�*�6����|�u�cJۧ��8�w���zuavEʝ��� &�M"_�S�������O����+m���S]���7q4�G�����(�k?N�E�T�RcK��'&�\��3�ѷ�y��JVe��z1쵣��x���ܥ��E���0KS�uA�G���}h��Mi�0��AOF��@�]�Gk��K;���7' �"��,�s�U�Y��R��Hv�I�>�H���^]E���iG4)�K�U��E:2>׬��1�c��u�m�q�ՠ.����?�fN~���F`���b����}y��������r�J���9i�6^r��\��q�D��5Ƃ���*�uy�5�$eY��|��ɑ����i\O��9.��1������gu���'/Tf�%�|'�S?^��D�I���FBk��6���z{�D�������%����-�\��-Ѡ�������pۤ�U�dA�C���!8�C���IEi ��vϘ�;��~��ɂn�9�뻭|&��IQӐ�]����Cv沺t���\F{�d�����_�B�os��i�׬V!��+].
t�n�ֿ����������|��<WS�{|�H��	g�*��]/�&��b�V�Nf�U���24���.�*��̺�Ҕ�B���B��y���`�8�S��\�?���\�@���x���Dy�����{85�ʬGi>f�ZL>N��F�-�֩���~*ضps���-J�4%�g�7��S/��=%k�h@^�#wh���nm�*$&�/��wg�������[٥d\��)a����q��yn=���Z�@aDܙ����O��nD����,[-m�P��{���yh��d�oz?=ַ�X;<vr��쀒~)�Њ|�}�r�q&�g�o�mH7�\d�K�>nk�AWe�|8<Y�i��Ay�p9<���ă�+��U�Ԝ�����v{TH'��%C�in���"~�L]���>\=������1H1��BO޷����FA̱���>-�|:]Bi��=՜I�]j��G��d��J�lp��g�G��2�c@x��v��T݁��u� s����/��m#*�uC��z�/�~}�1Ҍ���W�J�������V����t�St_Z�[U���E��%�u���d N��T�]i4����u:����޼ܿ���|BQ3`t�B�x�[�"��A;!�b2Q��b<)mn���Q_o�K�GŻ�.��3���5
ҹ�@K�5L�D1�7����R�����g������Ak>���Q{杬� ���Ա�4jx+��G���64�F������]
��O

@2�Yz�ʔW��8MGr��^�F�q�Z��7"%I?��1�!�(����E�'A$l��	:<�\�P�7*T����p4�������Ӌ݈�̊C�do��-[��|�T�����S�����)�4&�m��A���\��$��I����䴏���l\lUtWg|��c�@?KM��kQ����fٲzw����ur�MpPX�D͒��w ^��1�ƺ��ˌ�!%2sN��}Qx�K`VjjZ�o�
�&�cχH�Tl5`�BN��t]���<��p�����G��m�/������^�e�^�PI�($�l��k��h��̈́��y?y�@���w��Ӗ�o�!Z�"�/���\�l'�6T�Ǻ�w��B�pU�&��3�6��&�[/��K�4�YN�+�]L4�f5v���<zH"����5�o�Z�6�pH��S��SH]	3�t�p�в�x��D?w��G\�<M3�����\I�^�&��-��f���;2p_�~Ӯf�KIt`��|�b0�����G�1e�!����u��r��ap�+gY�F'�n�cŊ���,n�ί*���_0�r���y�֯,'��E2�����=���Z�l����Z��N��)� ����5��m:]d���>b�uI���' �xV)Lp�r�`��%�I�}�a�MtVp~�@@���'L)��\.m�_�|��y�����.Dbz/�I\0y���Nn��y�v�o}�r͵�0�=7W�K�,w�@9� �5cl6�n����v�p�J�jd7e� �&e�T�K­i)�|HP���s�"��k&䔢\*��f,&�.���gYO�����p�%6��B���Hy��uI��K�3�4��R�$(�Y)2<��P3������k����P�p �6����1��v:� wA�U2�w_���.��:FW� �<�xOO��D΢���c�� �qJ�p(fǁ�}bU]r�R�����}he�v�6S�ׂ��@w_��UC�7�Ahn�7��2ȆL8%��G�V
*��H$��F�Ƅ�()�i��"=�*�`v������b+^4�ש�:t`�J�QG�q��DQ����0di�5%uH�e���
q+��q��@&q�@r����.���R��w�G[��C��x�$z��MR���<
�֖�e�/ /������mh�7���S3D��h1��:1�V�A I��_���5��/�d���/�
����M=��r�4`�(|�>���7�}�s.�0�k���Da��|]w��.ʣ�+G`�o^߉(�D�⺦����&�p\P�Yު'^!���ƾ�WCE�����a�Ϻ��`q�[Mˍ)x���?���:�}g����W'�����m:FBQ��l�Uji�;R�P��d�s��t�1Z�T���Z��\���e����*v:�|�N�P���K�jD�i�P��50�b#֫rnޡ�����5lP'����#���F:�j΢�TM�3U�XX��jP�@X���$�\%��;��x��hee�F��ϋ?#���)y����`,�]��6�ư�O*V�l��*pnA��ښ����f�hhK'#� �U��>k܄��.�i�u>��8"��n�5�C�p�?5aFG�ٵ�F�"τt43�*���Y
�4�s�gI�@k��x�3�vu+A��)Q9u޼�[^fq����TI��Mkv9��c�Dl�+Ec�����@��\f;O�E�B�(��nRc�C�5]"V#��̸OE}��u�!�T���q�h�AbeIϗ�Ȏ��z��#8*��w��C���n|�!�sZ������*��o���{�5e$U�b�*�9[+�D%��^��Q���H��d�1� _�]�?�<2e�i&]����U�1�~�z��y���"���������<������4���E���@�Uk�E���`y�I3���2�$ČM{�����fD���P�ل��u�����Ϗ�<�}�~�ԑ�������s��s�ģ.8-.g8�^�.w�⽗:���cT��@�9瘯����y��75T��Yx߇ԑeC��.M��V��#3�S�6>(2z3�s�
�PC�푝#)��)��d9�@+~��D�m��\���I�]V�'����d��A�u԰��mt�p������l�ts"��B��O��^�Q9��~S�	��W�U��GOp���f��߯�;[k�e�X�?iP�.��������Y0>P<Ч�}I���Z�����h�y�12E+��FW�	��g�X!"*J?�SM���މ/��bvSC��%����Pp���~l��KJ�ʕ�2sQ�{G~nNN�׺������S�9<.�d��m���D�w��y�x�8?1'�%��xY {`S���o7���6AE|���J��A#	q?D5l�������N�Ě3:M��� _�^'����J����x#75����]��A�֌�޼)�x��������+�=k+~sW�������֟������5m��+��k�Q����C�fw/�1˵	0*��xS�M��a}ǧ��Wz�]���}ʃU�q|��<g�Z�p�E��y=Kd�8��>���.��Z��fv0�\A:�uX��!h;u6l-)�f5��CC�}���%�N:u���p�5�,����ޥÔ�w�^��W��ؼA�3�m�k�V��C�0�m43�2�Hf*i�/Ž�E�4�*Ӿ�%���l.,�����j1� 
IL�8��J�gU�Y*��a��ȳ�q֬b���%d�9�US.h��-ߥ�oϐ�(J���,�$��|��H���H�8�Wz���^J�dz��7�p����aWD,+��>)dۻ=��1�eo|�P��p^�fv���yxr�:��=���9Qz�LM��,������g}</�(q��U�RY��Uރ��j�+I]�Dې�.^S��-K]i,tc�'��\�]��-����<6xo:�|P��BWg��a��gUv`��g�E `�;ǁ=�<���X���|J����5��G������q�褤�R��/8O�cۺp��3|ф�̛�>��?�.�Uu��)��)�:���o��k�5�/��h��&������?���?5r��d�,�ᵚ�	���7�un8N$z�Bט
�6�+%��~k�������6M#����@iTP���V[R��s�dm�[�*%�����*t���L�z �:IS����X֜�������-A=6�]a����OWhv���X��j�D��z ��ή�W���F�X���t?������=���\��uN,�j�e��ı��.�/���%  PWQ����C)XF�P��񒩐�6���lk��g��ľGw�K��6�����O�q���|#0�'a.����z�kˁl>L_�����U+Z�,G��Sa�aHߛwo2�sejj��w�/��P�����c���a��(�f9x�w�������_@	
�[�ћIp&���(��+߆b4)o���$0�w�~ai��� ��N���Me��4s+1b��h;�ބ�H/���n��6�/��:�yR� >-K����_Š=|���ނr���7Q�)�1|WUdC��䚌B��(�ϡ�����$V��qp��,8v�#��~h��3+���v��'��[���>�MU)lb�k��{v��T�R�����2ې�O)1�Z���-ې�%NѰG��.8U�Z����W֧�R��U!l�E	��#ږ��/@�It�,�ľI���K�6�|�#��V
�\�Z\�Yj\܈a��Ԣ�*ˍ�6�|�N\#؅%�o~8��>�&�4�RZ~j�9�}9����3��ڂ+s� ��C`됡�R��q�I����0�C`����mtՂ��**T%�]�����.��7�--�p��Nx
D^7�����>�����[��O�_k�nT���<�As�I#��H�c�)P�$kf=�j��ڐ���
]q�#�R	��H�~K�/���$ŮQ��ܪw8P@�9�͞�#�S���\E�B���߮�Ts]���z��#6$�-^:�1�/#�����I�Q�mb�����Yχ'�%��j�M�mOp�g��>w�Nw��BxO)aSܳ���Z��)�!�+-ĢM��6��E4�I�4GUw܂v1?QQq&�j��"x%��G��>5�븀��ғ��ȉ�d�W��d�F~�!�����$b�
����[�{��- C�:8�Tj�ʔ*��bP͙8-�8E�s�=��ŗ��ݶ] ���@.@�1���H����䐫B7�������"dQ��J��<�ػ�3OGr��-3��l9a�ݏ��.��� X�/�>S���(���v��<�'��|��"p� *�)����J���.
�tH��~�V��!U'}7�smB0��}k�:6���γ�g��n��������>�B�7�u�p���)Z��7�Ǩ���{Z��+��o��ı�7�EGFN� �񆔩��J�fF��J����Y��ٌǍ�i�܇
���{�)ī������B8�wM�`=��2V����y�P�D���$�y>s������ǒ!H���d���F���.�� و�b��2��5�-�����d�S6N�f���,��e�'����6%qPMR0ʿ�MR�}5* ;�m�F� �2d[���Z:vW������?X*��ȩ�ܱi9��u��E;7_�����	b�/�����1B�Q����Ԫ�����	�],7� �5�r�J��B�,�D`5m�K?,[�(�ϛ6���g#[����Vb�YCp��#���P`n2������I��2��J������@<$��l�*�/e�kDN��ʗ�b���U(Bz7����T���A�s��~st��~)j축��@m;����*EIG��N	"�گ$@vw�+�-�
>RU��/�]U���C2&���AqG�I$H�	_۷/"�i�+T>��|,��R�KTAQ%4vNd �)fd�շ:��ҁ%r�kY|��B+s[ |��+�"��d�IjZ�<�Y�"�0v�	�L6��x�����<ǣK�&���[A��K���J��z�ڃ��+�$�`�׮Ͼg�ߑ[���Ć�4��ҷf|X�g��#d��t_`oIfR����X���D�������eK>��A�X&���A�I��B��څ�x���G�k���<=6,$V3t�����|�q$��?3	>R�ߡ�sK�?l� +S����d�y�N,�����5��_e:�y>���&ڧ6Z'mD�v�#�@qLE}P�ݤl�ڜG�eZ�PS��(6>��Ѿ���i򈈷�7�&5d���"c�89��X[��#8���-����j�ڏYx�E�1���@�u1�(��.q���;��P/�����+���m����3�g�Wea�������i\�[p���4.�ݽq�x���2�Ԫ���~έ���[Z:�7i}n"�ćRj�՜{A)�e)��,N�>�7��X��V����)�y�^������gH?q�;]78�D�(�,[\uEn�8OsLC}��l�����Y�#����'L��4��{�U�y�&6iأ�D�s1�b�f�V̬,�fiV���{�V"�E	�]%�U����[�:ZI�qr���'Vi`�� �����]�!��h�}b����3��{'!


��?ES,--��Cǂ,C�O��9%C"#�&Y��^?�,�'���*�g�57k��v�fO3 ML�w����T�l`c3C1o�sQr���md������-��w�P1Rh:���|)CR
�Z%l�Z�c:�d�\��&*�����$8���Yc'�c~�t� �-r�D�c�b���FH�\�3�_Wf�.�?4"�eǍ��w��pyY����r �$�}
��t0�����q �D&�
�]�U�\~�^/AH��� .�s�A���i6��nv>@���`�ԍ��U�������B �����5�ss�hy  ,�i���J��6M�MH~v�f�����'H>=��ɐ-��?�IX�a�N�Zg�i���˄���Ihj�Py2�̧��l���^My"��j��s}M�g��-��(e4l+���*F�����X�"��[YxK
�+
*{��+�J�#��^������UW�&cR3��bZ}4��܍0��x���'���'C͙9")��7��s"1E{��(�a�BQS*4�қ} �	�x�)�V:p:���"{�� �s�A�D��kYM@۪��g�z;̑a���>�ޝr�=�x���ˆ^E>�a�s�~���}��h��q�n��o�-����W-%�k�=�� ����Tr���-�]D4/�M��ѬN�� ����~��]���x8�f�������R�e�z���z�cY���hG�v����~���(\�
Ǟ��T�*j2~vN�xbH<|� �vCl���r�¿i��-H�,W�:<-����"Q�W�Aiéɩr
)U�8[�j`�LsS�G����_H�JW��.���\g"�?��8Fg00�%��5ԉ3R�笹�����<��w�3vVu?��-���|W�aYC"+rfVe0J��n^d��Ee:s����(W|t�U1S������t|�@1��]�U@��S�0�AT���p���c�ڶ�T��� '!h�f�����ѫ3/P�t7��>�����N����Z7��)�uX=��j��٤�b�6���f�9'ey��Rb/��j�u+��́�4���kZI��3�bz��.�L��lZudE��gvZ\5�bRq$Z���L�&ΟB4��Y$�����V~�N��鳑�9N66�`��/3��������AE*.+���;r&q�q���]v�� ؉��MX�"/ ��Ʈg)�� n^4L�d��.��n����,�Z�Z���-ͼ����@��,@�� �C��Nl"By� m�\�ƿ�u��,���S{��>?�v�P�f��`��!����%��f�~�c&������!�x��Ɋm���G�iq{�c08u��ōq&����!<���7 ��U�<�ƛ#������IX^�۟Em0��"?o���mvx(�-UP�����*
I;�nz�Nd��H�v2�����0��>�D֌��Q�쳏�e���ϒ�"�;����K�Y��ç����	��	���'�Xxp�,�S�,-3�-:W�a�ǢY4z����7<-�	�� Rfl�L_�_�����-'���#���Iv�Q]��T�k���9�H����YI�������j�}"��<��@�Tc����J-b5��Ҧ��aj��q�cp!�D�d��xw�v(0�Ǐ�|K"�BD�Y;4D"C8�/���v��M����;�ung��R˅(���(��6�|ʭ�<�sr�h��[+�d�����٫��KHM�6�V�]�����[yk�,R�7R�/���h�驽���1|�{M/MjgVX�1|[�<|^�Ȃ d�ew������h�ި�B��>���U����b�hk��#�&�����q�{����ԱQ�� �@$��d�2�a�y��U5�k@��.�m<j�;�4e��f���Q~����m�A��l���8�lti��/�T��(�p���oy��OU���+��#�m��^�������>9��\��(x*S�n���\p/NN���+]2������
�5B���������N�#���WV���T{�4��]�+���!Ř��B�����w��%����-o!�S�� E&+r�����VW֔]�w��0�u�a��MI��^}]��Z�8>��6²��$)�`c�=�.c����M��1(�/�xJ"�k=;3��Uũ�W��-��,#��?���4e�J7�W�����$�aǛ N�3�Ҿ�[�T8�L���q�q}��z��;��o]�~!s�D�h�2
��`�V��)�9i(����M�����!B���-o�w��?zd8��/pc�9�in�[�t�i�� �bp��Ht��Bm�@_�K�FN˨J�Z�@*�B�MWDa�f������tyM��UJ6�S��ŗuHv���iu��#j�D��}��~�}�j}:ۜ�g�r8�a�sv�ֿ���gI�4>��s�� Wa�y	�N�l���sdo��?հ��2�1��M�I�2ǧ{���\C�* �t��l"u��Ғ����MM�M��K-_������.i��
�����x�f�|n�_��>:��3S��V�*b-Ngp���x����Mg���qN˞�y>؀��H~3pz)�kG�����P�8�����qG��BZ��2�>jP�h�9��ǒ�u�ƙ��o��lssuQe�A`�)B�Y��ҡ=䗛�*��Wt�w�luOιM���s���I��wJΒX�>5{��`X�ps��8��nW�		]��^���(��l���&��R��3L�Q��U�ojH#�*��8�|�q,EŸe'.=��j���C�E��+��ߓSM��J�5n�J������ș�E���ߊ��A)�;�dnP^S3/�de!���=	�-�/���Y�Z�����B�3q����S�i��ёcy���z0"Ƣ�My��k�W=7�FN���Ħ&����U�2�{ �zB�L���J��m��m��f]�lk�iZe���P���i�Ž�k�<���a*��h�����j���e���\ɵк��d~~.a������E����й8?�<�=��;�pQ�o
\��F�m��e2u?�0�ij�!��*D+�ᢟ�����	�>\���qX��"���RCKS��*�"g���	7���y>����w��H�i��i*k���JUk�Qe�g�1sU7�r�XC����3\���U?�lin EI�U�j�|�Jv����=� ��«4�O�|�\\k�-�~yr��N�]{������L��^Z��>���>��g�A����b��GNW[M��vc�]�d��#��E���b����WPuT ���g��n��"�q/بW�ס��|�X�|
+/�����ǝ2Rz��_��tSGK�qI�
s�>���wR��pV�}Y�4��qqc�3��nC����|žL��	5�I�r����	�rL��s��a+	7ו2M��^WSw�0R����q��9��mj`�d���r�s9���3�WYX��[Zƺ�����X��X��p�C���#b�T����Mx�~"��[,�&&�N�N���F>a]$��3sk��5��y���J�J��+ܪ�:���	�I�+�N�b>�Uo�v/��h�a
�̀�g�R�������.?�tĭ�ҙ���?n�~����ĠS���g\	����P����5W��|���[����<�uY�6mv�:�7�fY���/wwW�'� �e����g.�gk�3�{�P�S��ht�B)��ϭ���\"o���6R,�-û!B^���U�&����X�GD�*�ڥ*�B���@БV���d���fL3i\�߰Q�Hn�9��Z�����N
ɕ8��SR ����Uc&��`�Q�'	~��h��au�! �}�c��S}��-��P(��y-I���0�X�����A��XB�ז��|���t�i�<���7�eƷ�W�Ih�z��)�V�3��2-��8�#T$mX�����~;3ѷ8��e4�|�kv�C�������54����s�O�G�� ���μg�#m.��,|{���oh���W�h9]�!m��^K_TS+�s�\�����vް�Z�49iq`��K8L�Һ�-��Y���.�S4B� s���[WIC�CsT&�h��qĀ��X9Kh�����w�ǃ�P�J��a�1��3%�!�a@ӳ���h��]_���|h�\ށ$��jt8��P*V����_���vn#ӑ]�3O��{c{.�p��ǟg,�Q��T�q:@t^�Oc�O��dƷ"�Y�td��ĥ(�6��~2���<}�Ȓ��)ՙ�|��c�[4�X,��s9�[�t�f��zo?�?�����{�~u�ٯ���Qp��6(�:��u���ӟ�2���l�[ݙ䔆�a��Ij�>q�U�Z��mX6�Ɯ�<��uz�:q	bay��U�(��((���(Xi�4i���3ܳ�
)I7�}��<��4HW���h��w��.i	)=�����X@C��
�Ks�1V��ߡ*���2c�����-�|yu��{�p� h��sxƂ��k��+-'�
D���w{_G���5(7t��1tzY7# ����4[ul��"r��e��i���SD[���U5dx�!?/-C�΄r�HPuUCt��H���b�������R��=���d���}���gK��P������zص7`n���O�Gթ���ʃAP�r����PU�!Z]��i���o��X�؛���h�f��$g�t}���\YRR��Z�ۥzw?�����О��NZ5#�*(C6yȩ�^�H"w<Kw�G����a�w��!�E��ݒ��[���!]^q�?o?�{��7
�m�2�5�D�Ydn�b�Y�%M�v�:��y��d��'x��ؽF��U������q(b��[��\�4J�vS��Ր��S���gwfq��b������J�l)�l�M�jm�{]/w��i��e��B�i�9O����&�Bm���!�C�������TVb���o��Y )$��� k�켝���f���v7L���EC�N����ֲ	�KZ��5a�`�[�X��%��0N�#�7���"Ը�6
�м�Ō%^�O�OC�?�;�,�D�s�$\��_�x��ܾ!�',x@�.�0������'�t�j���铂�������H�����SzS�;^ȅ�:,��|>��O����UJR��*�li����)�fx�>����c��������a�Gs���i#uZf������Dgo#tK)W�t�ͤ�t�PM�������At;�?/T��ڮ����k�����N�S���,��\~��ˍ�M�:9�I�w{��Y����Ód&���G Xt?����H�����}�/8ُ�o����v�ĩ%S���"�1�#)��F���ұ���(���4�*b�ӵ��f!��&�� /��S��s#���n��䩙pnii����*ߣ5D��
��ǒ,��l��w���fdfd�V��n�_
�\���=^��8��`Z�_���%��5���/�����>(d���4�E�I�ei]H�N����a��U���%ꖯ�[��*w/�'������K������@����պ͢k�z�E�T�GFcxm�٦>��uOk{��C�+~���I��
uH"AX:�;WgVLP�>�θ���A�=Ў���!�ʮ���\׌(�9#����C�&�~V2F�<�bL�_��#б�6}����<Et���~/MD����6�(����E��iu󩵎a�s1���=��S<�m0?�u��פ@��U�Ե���l�M�ȗ�k�S��~^2bi���f���W��2�x���~�+!<ߊ�B�z��O�8���?�!���+Z���v�Y�Lϱ�f�����w��Um-%���(��o�@i�:ʓ�a,5��Ӵ��Aa��q8�������|�'�^7]b>�����L/,'C��y��娪���h~�s��?6C��'I��_FFqM}�ގ�sG��?���x!,O�C�{D %����}ގ`��K.�D;}47����������:��>��|�ƽ@)y�,(�t�ɐ�ٱ� �`3�Y�_���3N=�Pb�.3"�>�O(M5��~|B����+����e+����(Z
d���*��o-��#�T��ф9�Iy&�}~���]9d�< �0���򅇊�����,��g�<v��i���Ч��>�a�jK>�יti�Le�/25*5e�%��4�
G��`|�z�Х�]����*�}J�!��/��<k�yI6Ͳ�]����!���K�Ƕ��5�_��풏''�qY��N'�&}S@ �Q6�u�B� ��T��;Z!d����D����A�5�,�|�[@�Q��d����+��xL����o���o,��vfޒ��A�=Ok��GϽ��^9�:p����y=��aT�h�VH��$9�;����L�'��\z�� �Ma����Vk����W1���H}�v%��/�WDI(樏���*�_-�)}m���Xߞ�z|�o����F'��>B�/=ncN6x����V����888l.�@S��[��Ԣ����`�����[���>�V�tKr/��i����I���΍D�i;U#�
���릞0ѢY���:�$��5ƕ�kÒ��!��ߐo��Ͱd�`��f�_b�EAm����T�ep�A^����P�7%�S� ���q���#?�'���@�
���S��Gbi����!J�V��){����=�fbf&�F�\�3x��`P�A6���q�Q��>��J�X6�!v�M�GL���m.6M;x;�͗{�99-تe��mP

�E0
�H&H�I}W �zNX��hm�w&���}۵���;Y��l�J�+�&Њ��o��z�E��5���ux�S1-b[�JW�}����Zm0߭j��������#�����6��F�^9�4>�j1�i63�ų��w<ХX rfxż��^譪��m�(���g͗m���f�~�����/0	�%��D�$��&v���`k���˾�Z"`:� �'��40aNd^|��4��l�!�r�-Z�w�A�+�l��4.��H�����>�Z@��_�S�f�w��u�u������_l�|����`��R<'}�c덆m:M�c��'A����`�����;���y֔~��?�v��(A������G�O�+l9�5�B�o�$�>�|>_�<ȉ�A�cgqt��bV���� {��S���ۺ>�,���B�̾C��c�fp���Uv����ՋT����u��N�Z;�������~�^�{9ns��=�|��?$A�F����R���c#jo��ɹ0M�!�?��.�\�9b*��W�?��`����|���v�\9��b~�b�s�����\ܐYC&�$i�Xǭ�����eZ��̵דJ�Eҷ��͍*k<�Xئ5�&�C�1���	2�_b�lT[��?�}7������n�v��z⟯�ػ�}/��U����<H�v����8�se�x޲����_=ܟ�Jhi?�`#�DL����0���0R�Mx-Z�q;8��Y�G�&����d��0�R�i�B*Vf�����p�#<3:������
ޏ\����#�?I��~�%Md
�M7'���[���v~G�_���CΘ&��,f�2{$}�uJ�O�%0i��,S�F/��W6y��C����IL���_L�������A�SdJy~�B��&bRA�ٺxl(O����1���3�?6�e��0�����D�>_��c|r~Z��{�����r��o��BϊD�0��Cc9� ���&�n� ��D(AѸ�b�;k���YD3C�m=��3��4�XO�Z<"������@�mPi�f��Y���gZ�� u�D�G��){.}F�S/��ٿ�ت~�V:���0�����]��x>QI�#�{����w#^�w��u,���ò,P�VE�X�o�)�#KU~��}�-V{�\�%�vs�N�aEYB�4��M�PL�M��A�8�v��~gQ��S��%��Z���A�o���ajDǞE"�23�R�q����U�i'|�����������$�w�0��:��dSx7q�J�5�������c)Y_s%e��4MR`���&<$��EL�'�/����H+d(�Q�_FE����r6肀�Q�.R9�6����u��!������_l*U�	=M�$��#�K�M�>����M5��@�掃P����j�U�/��L�u�k��%�4�S�?8a��l�f.�gnc�׺I�e�*��+ArYH*��@�ú�-�)��D�P����Qn�~a~���P���l�
Ј�I��V���i�<��2����eP�h�SQ��k���ڕ�K���E��@kmr��r��%ZNm�@��aiB����D�����Jwqq������_��b���D�S�'jD��lZ��m"0P��`L�y��(Ĵ��Sė�?{�86��ϯ��K&Y�~1��שB�4{�k�{���:S� �q?^�:A��p�z�Ŏ�&_hn�mh�գWS�d"�'"��zV?+����B�x;YY,tc�J�ʭ-�(����@���8/�m�	픈B\�&�qo8�� p���� #<V:&+ ;�Qf��t�f0qI��Q?�����K4��Pz���$���6�^�>�$� .V�X��o����;D�;(`sm�9;<|(���e�#�,�ߟ"am_>yb�A���D2�	ļ����j�$K�,pd�9�]0,'�J]U����>v� Jh��s3��K���f�g׌�tI�̞�"���y��^|{zӨc*�<�(�s ����4�����)1F`N���S~L��O�+?<:��Ef&qu��Vlԉ?N�;9��E�&�C�$+��2�-P	}�Q@c��R�����u�	<����0o��c��_#��!dD<X[�]�^"�7!�����6C�Q6f�89�Q�Cx�C:�Z�ӣG�3-���P��Q�JWߙ�O�ْ*I>l`2�z2������A?=b8ر���ť�C��Z�.Z8��tm�A�����ja��_�GxӜ�u]jt
<^G�T���&W�j#b~��=F�1�Np�{j)����E4��I��o2���Uч<�	�����g��ϒ��5���t��?P������.d�������6`�"D� SpZoa�I�N����ʬs�ʓ��x����r�O4	%q�L�����ɍX�0J�1<�b����<���Ñ��on�	�]	���­��lu�cG��/Z�xd$�Smu�JYP�O 
���WE[���/�W ��(tωg��bÖ�K'�7q(���%��)����jT��̙6Œ<�Iw���)��(����o�{��-���'��W�>��a4zj�X�6TA���@v�A6�*iu`�p}�e��˚�x�y��#ѣP{��|(�τ6ZkD���
�*��-0~mWᲆn4���=�a������*�)��~���֩_U1�q7}y'���H\�V�i��x��Q�E������dKAJ,׌��Xg��x��2]��zæ#I�qK�=F}��_�����_��↦���d�s���G�YN�A>��qli3r�&E�~}��]"S)e(� �~�U6�bߢfv���W�è��|��QL��k�v!;T�Ey�,E$5�g�\�j������[f��f�i�v�0d�mG�3����cu�0s��2u���[E���o��G*{'�f�M�2+�^�|hL�4�K����I�19�(k:P�B��+�̞�M��gEF���Q�v�bD�P,�!�Ð>c�N�I�{�U�=|�}<���`&�Kt8��
)���� t���eI��B�*�R���XJv#Z�;��w�ԛ���W�Xa$Tn�5;w8�{�ŷ�-H(����q�V22�:�`j��M��C�?Q��Ν\��BRޱw��Ot4��B�f������;¦���T.[XS63'K �*��N>KZ�Rr�����Z��oX^7����\��ط�a���?G���ܿ�|@�������Mm-8�Yp ��U}Ӆ�8e�� �;�FRN�5�}*����1�nOa��!�� rq�X��&�D֗��Z ��wЦ'Y��dn�o�RkPx :\?�r�2vd��'f���W��R2,]�R��'g��7'"��{*�a�2�O8@�h�>1{�� n���M�Y���A�rnT=�K6Zo���Iq�U��9�"��3����A Q!�&B�0�:�!�ر.X'G2��Mc�k��P�������7�����F>|29�X
9�N���@>�3B�.*�N�������X���������ڭ�����(!��&8��n�"A�-ݑy˒\Gp�udeQ�oH�1�v|�e�3���2Q���:7 �ދ������~����4-.Qu��<�<6��/c��877�=) d��/��r�b�h4�?f�X��7g���t��_�j�ۂ/;�B�AY�\�j���� /�����#�rR%3�VB�.�ol���T#Zh����GVY�J�<_>f���G(�K}W�bts(�+4�ğ��Iڠk�{�*�h���M-RЕM������:��6�ҿ+�S�*�Q愧bZ�;�m�;M�����A%��Wr�7!�#X�Q����ծ_���8(�Q�Ѹ/�{��x�� - �,��z@/Bp����<��"��j_g~�T�tTR�wS�>�p�>{���J�8��?��R�c%
��DpsԆ��&�qE:�S]%χm� 嚄Ā�8#%���Ւ�f�*����'햵�|ޭ'h��<��
i�\KC�Ǟ>�*�sM_�_a$�@tm�&9�f�����G�	;�����}M������(�?��e>�>� ���[�_L��J��iFw�_�H�:{=�k�{�Sn����s����^~Y�weu��Z��}�1./{Bǽ�� ���m�`�uj��R<� _�J!=[��n���jD<�e'�- [T������mSRr�R��&��"��z�
�Pڲ�>��H��q���K����E����֐���Pm���z'n��q��ժ׀��m@�UOS�"#;�#SM׽�C���!����=�/�z	���@U�����`�>*�n��6�7��6���x�ћB��oOES�yzr������ ���
dp(����U ۘ"5G�c�N�ߵU~}v�_ڿ����͉pW�0��b��\�P1�/X�B7�9���h
*�)"S�o�{�mz[��T���}�08�0X�o�q .}��r���p���t�`˿�?�ҝw�L^���S��e�q�:�X��v���n�o�N�褗�����rz'!To!�4-�#���N��ܔ"�c���]�;�:Ԕ���v����>WS�i�B:��6�q�	 ?5>ȡVft8&ӴS��2�A��ǆ4��{��N'��Ʉ��~N|�]P�T!�o�r�u��#,jRȃ��)��e�U6�7Ç��6j�㫋?rL5CD�^�Lo�??mE�`h�*�x��i �֐X�ص��Zw�v�+� �Ur͑��=S�^]�tޣ|&��9[��!�L���t�H�N�:�,^jI[�l�_\×o��������o�u�[���r4�m Ys��>�|��q�*����u��DA��p�\��-���N,��%f�����1'Ջ��4�lg�3���q��V��;��f�9=G�"o��?�
B�+}ӆ�m��P�~���i4�"�XG�=�X����߿�$��s�}װ7(H�X�t�N�w/;e �S�gmox�2��c�ƚ?�2-�R�*�@��^K�r�(�6&qu�GƈU����u[��x�p������$�"����%�+M��sh��-Z�/�����@��� �
��+�٣'�.�S�\��M���/{��gm�L�)Ԙo~��j���gQ[^G�|#�H�0�w1h��U�S�sBJH�#R��ݴq��O��]�c˵Ʈ�Zr�����]���G盎�v�-��)˂j��ͻ��{)�`x��e��HU�-}������Buk����C!�W	kV���Gf�i��n�MM�=?�+�b�k��B �%�Ol����{���u���K�v,���v[�ͯ���+? �<aOJ�Ppm�*`F)1���ľ�S���J��� ��Ĵr���\T�������{��9�n5�HsrP�Zt�X�v�a��l^I2����8��v�� ^�����j���el�'�m��0Z>��<Yh��8 r�������1\�L��I&S���9����&V�>[R�0��e)���N=�h�w%�װ���GD}A�Pr^ee)�r��l�{8FՌ܆�/��J���ԿMI]�;7ǃoD*����%�kX�[����X��6v9��;J�#���;���:�B��}$ ~F8K|捑H�X,|y�v(�zm_�u]'�^'@Cp��z1�˳�bN3_�9��:����MLW�g�pE��|ɾ}�c�/��k�K$��T�S ٪��|בS��V(|� �{��R�,(����!f$�儶T���\7n��r
�'4�^t�8�����O!o/��?(����=�
��r�
d�K;�{\����2�\�bi�W�nt�	>�RW>�J�u�}I˦�O��^�Z�7k�}�v�����}��PI��oC����.Z�O�[]�N2BV�4t8�WOs����β�����|@�5��g>�#*1�р3w��`�T�n>��X�u=�p���;q�{|(hT8���@;11b��gb���Q��� �I�8��D�����t,� �����m��Z-_&m�ÖisCVhǡ��/��@�U�q��X"�T�m���/��]S��=����3�vIGb؅�������k�^bp�oՉJ�U�n(Wj����z���p�|�{=c�����ģ��`�ٺ�@�A��D"F�󵧳Lz޾��\���x�!��ű��!�7�6�O�`t�]$�$A������_`ት$؆#]�h���5처~��$�`�@�]	�v��>�>q1�u�ԋA�wކ>爝_��C�EHF5��0�c[��Q�D��#��+�Ϳȅn�_��$��Ͱc�q���kM�<+�֙���`XV����ߚjV�n~U�v�Λ��|����:��-n�b�Jy���|tupxrI�l�_]>��b���
c�U��������BRZ;7�zBx=]dK��n;��s�k@�ʚޙF�\=�˶R�Dw��TC�'��M��V��a�+��T�E&������R��B9�\�Tx�kr�˗l0�� �C���#zsC�"�s�n�Ȯ�ӱD�r{�<o��i���MW�hxC���*��Z�H�/����׽�W���ŮD7e��Z�E��k�ڶι��Խ�$�ū��֋���=A�.ˉ1:%x�Ϋ-�e�(�r�E�%��i�y�s�>����#�+��a��
U6�YM ��ʭ��}�X��������^#憝t�^F�+����j�'���Tc/������&�`�̐����$���:�B�� țT1×ش���L�Q0�8ë�oО���Z�s�
�ߛ|�ۡʍJ�;ݞ���Ε8b���C�w��Qˀ��S0�����	��� ��a��6�QFȜ��@������7a���_V�];h��LZ� �V2d�}�ᅁZ�Wo��\�Vo׻?~���_c��`ނ5z�q_��OC)�����C�w���;��g`�Z��=�0�A��%�e��kC���S��c���ށ`�ƣySG"�`s����1&��	y�"pob^��� �����h� ۑ�_��D��� �7�ҧ�}W>���A,ڦ��pp8���G<o�Bnv�t��uU���Wɵ���a)�n��"[�?T=���X�*��zS�֡����bͬ�A3��O�� ȲϢ�#�t���8�7��7a��߼gO8U������T���wc��X䀟_�_j�wC��lE��5类/���mb������QPóÙh�^tF��+�'�7iH�<�����]�˥��^ri��J�!�ҍx�?U��+C�?ſf_� ��4-�d�r�����j�p��BZ�n�C+�TOV~�.�(��+�+��-�.I�cyV$!{O����5ԧhOײ��r����;��gc�'��㷙C���*&z+6q��������l9H�!cC�ځ�����Z��P��ۂ���Y}�ت%w7ŷ�|ikfi�1rܟ�#��(Á���A�.;-�(�0�r�+q]��x��S�1�Sp�-�� 7�!X��R����X�É�h��	���@e���A7{���Y��~�W�������T�(�+۝����t�	|f�%:S
���΀��6��o	~�)x�a&Nb�Q4]G,�#�$ۭ<FBd�s�3���Z1�A������wv�N�h��b�l}�)�V��=1>O�ɂ2�'��%��R��3q3
#5����@~t�@��|��U�L���T�Մ���km�>�?������S!������/�|4��A�������?*��L`�E1��CJ���2�Ǆ�|^��U�;��أ�����y��� �=k6I7�7��*�v����J���N�{r���q�V�^�4�}��b��~j�c�԰�o�F�p��x����6]aS-�͂��~�����ݴ4 �f[)얅ٿ�[�v;��s�kq���7�j�[b3CdæK�ח|���*х����($׷o�)q>QU-�I	��O���@�P1?Į���L�̲�q��ԙ(,��˙�B�w�H4|s��n��
>�B�\��8��y����"�kHMI`�VS��1���O�D�c�ئ������W*��U�Ҝz��$�iֱ������q,Q�>g:�݉�Y�:�}�|[^���.��Έ�`9��ڸb_�?���G�a_��ަ�4�����Ϭt��5�L~Wr�}���7��c��G~gK���~<$�"��%l{"m��� �o3�i�6���+�}�,B�i�L�«H~�L��Y_zr�3j��8^��͹�,V��~9�r�Z�
k��H��*��wZ2�\C7���Gj��/W����jL�lu��Ps��_���Kl�o��2S�����G/�w�`��op�=�jr]}����1Q��f�֤�YhD���-�Ʃ���A��ƨ|�;"�%^1e�ّ���r�������/��1�-g�g��U��i�h��9m��DBlv�����"
C�J�?�t��7�Nuq�������~̬�2-MS�``�d��|����L��F�͌i�'�QIĩmGBm������ܾ^}�5����f6]	�/�=J�����ߓ��0+םi罯��[K��|9��k5�!�k�e��1?�bM�'[�����~wܵ�U +9��"bø�-�!��Ŋ��� 5��a5lJ�լ�>j�b�9����5��D��s�l���w���M�l0�E�A���e�WB����|Egx���5>1���9�~���;oR{�J�=L%U�u���6�Ak�p�x_n�6�<ծ�Q��`�-U���Y���;�Ɵ�9'��0���3�����\��� x*��^Tm��(��£N7���3���Գ�q�Z���7��jb꣔��\kE�:�ވ`zc�Ejjn����9|��պ)����8�|�Ǖ��YR�$�Mqof��vm�����&�����ä1-}I��y���8$���"u��QII�y�:]6;@�$=���eZ����Pa�V����:�%�I����
�S��яW�}{��	%��vּk��g����=ÿ����"
���qR>������Y))��[ϼH�>V^����{�υ�6�����L�5oݟ�e�zlz�v\
ⶹL	ښe�p�(~�x�����H�a�]�,��u�Q���֞�͋�������&!:��xV�tn���l�%H "�I���������k�e!�R�sO῾�"��k<�.��[,o�����n���M�8�;�/���`��C������x�KHĚh�J�)%���x�F��r�3�ɠ��(""" E��{��ҫ�@轇z�""M$ z�5t���;�"Dj H�p��;e�u׺�_ɼ�wf���3��'+��T�滚w�)��>���>�Z��J�(p�%���.L~�SKl���hS-U�eMίK�_�/n��{���Ż�Xe�js��σ?���L���t�o�8f�ZO��(�����F�I���8�������#qךdt����xV�Qߩe��^�]3{�Y�b���#!���<���U�Ѕ�Y�=�7,����:�A(O,a6�X1����3p��&E�8(j��)u�z>e���Cdi�W
tm崀��ɻ�̉�d�I[������˝��%��ճ��^݇<�+�D�tvU ��0$�]���a�ƶv���՝��:�U��[]]�n2?��|$��!2.�p�����`o_�$�'m~�akI�ƾ�!%�K�"�E��m�������r��S����F�S[�������S�4σ�ƪ?��~�����.�L
0����t�>�5*��m�`8)4]6E��@_E�����]�2��WV)�4�7*�Ghf��+ZIw�|��?��r��q|yZ�W�~����3N���Hh���:*G��▥b�l>AS�f���yZ�̤�#������������J�f�<�I���9��Έ�u=7>W2�av�S�144d�TAf����'�Vb,���$�v{���:�"G"$�+,�0��ַ�N��G����%�Q�5�CJ�t�;�J��h?��a��i��)\��K� 8[y�fc��t�r,ul�=�8��_�U�hl�3+m+4'������<��c`A��N���́%��v���؅��s��'����ll�cz_��S��4
������w6�%H�����_,�O]�]��';���.۰��׬���@V`�W��>�0wU���"�m�N�D�x[����Zr9c7.ŏ���� Z����C4L7���7%�L��$�u�8\K�x.뫝W��V�����Em퇞L�v����n� k؆c���6u��#�_�Z��E�O�P�H�]��b*��Ϣ۝���ҵ��-Z�J{��0v۴�?i �t�dK~��ZD��Z�����<ndک[+�4�˴L>_m��7��L~�2���<Q޴=��߮[�PO�B�n�YW{�	q���ka��#�m<���� ZB��u��r�b����ehA�>v$ط��"�EB��W�nT[����o�j¸)�����xH�֘�7Y�X^�Mb��p��n�zԓsF��@0O����n�5�~��(��m�O��U�NT"�+S�;��pʟ���#�����0�h�F]����\�"١6Y�4�)A���	_,�����μ�m~ݝ�zT�
,�^����`���6�\Ǘ������X�7�c�M/��f��dQb������w0cb;!,���1ݸ#�cB>t��<7��N���d6�~F�ݼLɑa�EK�N����`����j�F�iჭ���gF���P�[:0]�Ѿ˚��Q��| �QqX�6�9���.�$����u�,Z����c9Fq�W�.$!WOMS0�|��oJإ^�b�jQ� "*Ɖ�\>�P԰�*5ϊ���e��F~r�6�:��g��5wE$��/�3}?�wt��������eǊ�AV/>�}�N;�CdS�g�"�WiI�}���T7�؟��5���E����T�����m��D��G�7ZM�pY5A��H����%G�\v�Yhu�^�9y�eF�g��_��s��F:��_E�@��m;�
��aV1#8D_c�(-7���Y��Kba���xpB�晽��nd�[7R�0f:;ö�[�y�TMZ�/	.\ZPs:��*������L�3� ��u �"o�X,�#7X��	8A�o�[�&��A����ӱ�/+O>SӀ�D��n���6�![��	2*B�Y�zrPBޔ�j@���g�b՜�����($�r�9ށS�sw 0Б�Bޯj�.�U�@2g����ذb�3.#�,#" R�$�4��t�F��jdH�9*V֪����1�A�������HM(�f˴�ˮT'"!�c9DG�o��a&��}y� E�/yn9T/v]R��2eU��GE���b�"cG�x>���p�A���%b.��Y��p�$�'���`��]v�,�¯n,�'t��+}ڒ�R(u�� �ȣ���,$&��׳����
�F�|�L ��'�".P�$���O|�x8���i��BV����*����q8�b��L���=G���Q�J���;������:-��B���0��c%�-�'6nyJ93;�R{����|�*@�o��/��>@��``��1�h�E2@���^����'�Z�Ƞ�v�J�}�~0�n�-{|��	f��sQ��:� ٞ�����a�R!*';R�^󜅥}*�v���Ier���X�:C�@�؟Lχ�d�����u^��|� pя���>��C�rp3]Y�nf����.�k�����f����>ov��U��x�'`j:8x,�[|�	Z	t� T��x��Av�JӏN�6�4�)�P�Eq���U���z1z��u��x�~&ɮj��B����Y~3p�w����*�z�*-�o,h<��r3fj{b��4TsE��>�1̊fh��U�=��pwl5!�<���͉9���|}Y��z�тNu*~&�#k"���O���3���j.��$�[:9�)�M�"��}�P�Z�in K?�n���Ɵ5��/y��_|��V�1���Ů-S��c���`�#UI���>�ކX̓�7��(�Cj�^��R��겡e��ȴ����7�����}/��ٿ "/Mϻ�b���g@��Rѣcp+�B��(�%Dɍ%?�']؁YM�4��y��:�̜�d����:�5�"N|X���P�?��b�?ɖ<���c*E��T\xPר�����:����h�����	}��K�R����mlQc�4ʇq���e+A�N�Ѥ�B	�>�#���{L�7�㘓��)@__��^L]�c�V̽�d�p;��}��|�pl�ſO�tj:4&�BS���Y![����=y�T��;�թ�xܲ㏝�/?�H�&:Aly��֒x������;ZS2�/J%�����'��-��Et_���H/����jxu���vZ}�Ώ�"ڄ��g�m]wJ�Y?8Jd5�5�Pݘ�Jy�T�A�C��	`��}��6Nޮ��+�NB�z�����C�濲�q]0ĳ �w%�t(��ǲ���ui�b��ߥΫ}��Xq�-]f�m�Y�fq���r]a������`}�������ڈ�� i>_�����}�h|�B�Aro�$����nu̼ې$��j�~N8 -���[K�Ij�RE�����2=�b��.��~�x}���oN��F�F��2ĩ-WY+R~&eU�Q��\I�9�o�n�W;Gu��`L��1���+�汻܋{�X�V���1�M>HM*M���v��T��$]��_�y�P��|��@��z�\���}[<h}�B�y��x͏�Qm�����w�%�&�Ї.,�D/:;��Z>9l���&�{us^�	��	7 �/��/�.�ͽ�&�>cx$����ávo,��s��|_���Xrq_�l�B�	�u
�@n9�w��
�j�s������V�+���xbB��%�s�6c>(+����W<��t�Ά�&�Wj�ĝ��S-y�f�ٗ�]����Ɍ˞��c��#��e���2�ɫ96�X- |*��ڥ��dP�+CJ�K�~��^�c,^�D��E�6.��<]1���>�������C��%b74�.�P��Ƨ�ƻ���;��0�cV��?��3-ח;�ȶ�6��F��/��X\�
�)��.�N��~ʔW<�jgΤ&��������JX�;Ôc.z��7�
}���w�N�X� }:h����	�Տ)v}ێ}δ���őixS-y�+=����Z2CB@i�&ݡ�����F��	c�q�T��?k�-�W��2𼧊o���ڻ��{�/��ɦ�y^���qq�s��8�Du�Q���3�ie�(�F��?׷^#��ӻkh��t���[D8�qT�)�
л�6B�uu�)�hbn�'m׬��J��,j��f>�Q�#j�)�c�⛵��^7�{��ȕ(��ت��]a��[�~����8%�c8�s���+��1ܣ���)Ày��}���C��	^��%�'�>?=z�F�4Az��p�A���s&�%f���Y7Ğ���#��6��4HC]��c/u�o����1�<��>ov$��ٸX�C���6V��)�*H�c��p���2Ó���4�a�-��9(wZ�5Sh�ܶ��/3�<E^6޲��N�5Ql�r�xգOJ��z��R�wS5���ш8��vVܶGh$T1����ޗ�}�%}�5oN�ۦ���\�_��F�ף��Ո�2%�Wժ��~!u�s���A�R6s�m�v;YmJ�~�s���a���◍���N�v|1S�79���7�i`_z]�a)6��4�rc|�s]h_$W��lJ�l�9�>���JuY�b/�/A��;5�>4����{bJ�Y%7��7j���zcA��5���v>�p��F�I9O��O�)�%Q��: 4u�7��ay��D��u�B�W�D<Ȇ�Ь�+��Ԏك��D���Q.O�]7�c7,�u�G�:-�����-[z6�n|�l�L�I���h��FI����^}3�]������p&��g'�&�%C���=�!�0��i1^�:���\3�?���i����G��;��١þ�i�=_5�
�����M�~%�8e6�c6
��ڹn5�7!��gf���8o�9��^<�?޲�F�Oy�'�b"��<�:ju��uN��W4��ˋc��Tx[�[N�y�Ԓ�pzCa���L�����"L�S�w��\�ބK�94��56�J>�P'�֘��y�@��@#`������ ��1�eMr�{�����6��?p��<|3�UWy�����(��7��-x�)�ֱh�v��������ה��Z%I�����6eP��p3͆k�:`���d�B�^'떙H��>3��n$L��S��^½�9Y�Cb�G��l(dGu�a�M
&�0�dn�rN�g�!�������K����}ѫ�$��[��9/��7���
y���F݇}B��'�����}�h�P ��F������R a�D偏V�U�?L��~2�w_t�Nz��^�OZ�C���,Q��:�$S���5�P������}�K]�TO �6`�:���5�L�,I�]آP�N&WNVy���j��3��C�>�ے�-�Ű�M� +2��\Y�P_����J.d��s�ժ�B߬���Z��:�}��B�8���SY�$.�eUۓ�8�<����
l�0j�	����m$�8��-�j~>��ܮ��|1�'����7ے�t�%�ԭp��:�T�j^>w9ڹ��IdV��6��i��uZ�A�"�~Ib-ˠ5}i�)���-�>ͪ���|�t}� C�|?|K.����]Xm ���:��r��_�����(�;]������~T�z�|^W��4{�M�W�ۼc���@0yz�
����N�7J�ѾCAQ��ӧ�������}r J�ۢNN
������(o0]��J�d�8��֥��|B�Ψ�j��c ���n~U]�ҽ���p���/#}�-��NR���ݐ ��䥧Z�A����+v��QH2gJ�l%�%��a�|!�R��p�H��F�o�A�/2�+��u�:��{�\�,���o�b
�ߺ8+�M"KΑ�RO[F����ͯQ�҆1��[~���')�TqV>Dg��*N�"Uϕ�9�A&{:����m�r�#<���dm�@Y{L㒕��Y�{��_#c��)�p�lfs���,"��"JC� <L��d��
<�(����Թ��/Yڧ>���|�!�
M��:�qbC0�vĭ�E���ީ��,�C���������@�D��Zm�����	u�dY�S��(̴� ��$1�G�+����<(⏭_��yFV�����t��M����m��s&��ҡ2�)�q]a}i���	.a�2�����w�RE�l�OC;�Tr����ǜX�oK$��U��������i����,�$/NoV��i���$��=Ob�V��R���c^�n��y�\x)��F�� ��j��;�#����?ы����*K���ἧoO�R�@�ӕ�a�O0O��Z��vQ6�iދ+�3����ڱ,�p��k��%���ӎ�L.A(�ck�f�J��,sk��gT�V戔�����.F�k��=0��Z����#�l����¢��a9����Ұ#XX�j ��q���u���0.�*`ߨ]YAV�0~6T/��À�S�[�.���*�:���IH�k%�� �L�R�)�p�o�֟M��jo���n��ԫ�;?߄r�'(;��cjcep�,o$��ȎX��8�;K��^����]�U�=!�)<ȏ�'4�ev�z˶��;�%c}��SB��"6�,�"�ݚ2e�N�"��܏�)z����<-e�w ��r���e�n�ܦ��O�I�2ϋ���a8VMǸX�L(�߮��s,q.eV�:�T��QW��gM/tq���jX��x��˭��TZ˭ ��<p��f�5���_~d_v�!7�A�� ����թ�G��P�R��w� ��智6G4��]�ְ{���������vzN�!��ݡ��ċV����K��BVB�d�H���L44��t,��-Β[;������h�)�-�����']#�CS�]L��-����yڞ���R��&��v�nM�/ݲG�����)J�(|��D(T�E%�Q�@�����w��YI����!.�<Pd��Sg�*��_q��mM�+�{ I45Ai�	��A�)Cj�RmY��8b���G�T&JXQ-�*(dn��^���K�2]��_D$W�*(%.�u|��P�/p�\ I������$�����7��W���pjG����@=!	��R�n~�E��#�F�CY���3�É�Axϔ'�^�_�+-�YRd5���\{�\�ٚ5�+�!�����iZ(gڄ-��3Uib����j(IqPe� C_,@v����)BU2Z�������ߤ��ӵ�}Gܼ�5���q}$��k�^�+Q+�W�6�Ą��F��b놔�j��k�{=91ð�˥�mϕڮ�蝯��#���駪��f �x�	��z�[8Sٸ��F̊_�f����`����6�4��"M+S����cq�� *��.]�����"f	���xq^xE�+;W�hWϭ/i������b���ݢY3['Z6�^j�nϷ
>��T������/��vw])�D����%Ie�ߪ�g��3%p:���k���ˉ�ȷ���$�_�$��������+&1�?�|G�X�����6�mF�D,��������.k&�7c���u)��yt��DG5��}Ь�c7�ͳ����w���)wW�N;Lx�R�fb���Y��-��믧�����wED�����������1��Z��$i@����Z�%j ���)y��!qA'�f�<ȕ�"g+�孳
���u�Tǖ+�l��D9�0�W�=�����ꩾ1V��*�[��'�z�۝����G����6n�Yu���+<'���f��D��}+w%�h�|. ���:��f�ɧSM?������=��8M��u�6'������)CCB�"U�������x4�<q����ry?�p6�p�Nh�0l�eZ��A��Ω�Òxf���Զ��v9��M�
s#k�S�2w��Pv��<P*����|���~������+���{�o���?��I��S<(q`�����B�Ȅ'�@MF��W�?sNu��ѧ��OeӇ���4L�݈�X��q�$)s���ʁ�I��&�K��a����ϧ:F޹��~`vA�P5��J��H5-�{��c��E�O��f���b���a�������uC᫱�gKL�x��s6�+v�"I��Ć\�>��/�%���75��*�� ����\X��*^��GC�An�F��&����7��B]���4Җh���sT�U86ґ��t�|Uٲs*6����)Gտ�&��d�A�hr1Zp3̑�_�n��8K��/����VK�����Sͧ���3�e�פ�'5�(_�Nl�k�{�y�|��7�u�&.��j�INk��=+�E��<�>��Q��UY����eu�Q՛��������<�MDPy|m�>7����3κDP; �������Z�t��O����3����u��'e��ʣ�
�i�{L,��I�c�hY���q�EUU���e�o��Ǵ�5�j!�N8J��hYto�P�D*_�[
Aa�F�/�?�,ĖPi����{���a1�I����! @�v��?��wXDF9ǔz�
�tV�_rb7!z}����>� J�F/�w�T�!������A��{�`�I��,�v�Q�ܥSUB��`� �!�;1����B�}�� ��Ĺ��i"F�pRKԟ�>jj
��it��^9�]�j( ��]���W��i#��wN��RuZ(s�ǥ��cvZrU���i��]_��"Q1��+�\EKR�nn�����c��#,LgFǍS�q���2�O�reU��z0���Ux�gh���[�4D3��k��; �y#�U���Ge��?������M�z�b��j2t�QS� t��W'�(b��̃N0֬�t�5e��Vf�t_\�ėC�4 d!k�vE�����j�NNO:����y�'=W�A��k�e螡[�-kw�{D�õ��]O��_s⬰��}�h�k�����)��/��z��QO�̗fu��i@/;~�7N�ϓ��Ch�k���˺��� . ��K����h\���R�@�M��M�j�~��7 )��5r_��y�T�\��Qͨ�)
���ԧ��چH�(�}B�JU* KL�l�16w1�0]�^Z�
�Wk��F�G��)�I�Y`1UE�jz ���\�Yk��ξy���X�E/-~�_٘�AU'+�Z�(+�˄5�=��'��lF>U��������P��Ѧq`����](�t����f�:� [���h��?#�oRy�v��7 `b�����g��r�(�k�6NNq��KF�f{������ߛ�d����@�i�+���GX^6�����6�����l��Dq[��CWV�����E/	���4ʷ M�|FKb#5�l�,�y���p9vǪ��;�j��V#���3dH!�R���=c*m�}ŭ�4��8�k\�cQY��_ϊO�_�� �`���Chq�?����*��՘�-v��=���7������s�b��ܮ��蓠.��S�7���'!]��~|����C��hdR��x?��aM�]��m�V��{�G&ꏣ`��A�"W��\ ���d��d����AX1[�_s6UU�n�7����M�@~������=�P��e�������XYHj{�r\�]����H��W�M�͖~j���w��_�j����yp0�K���"a�K�Aû���T�Îlq3�mf9��ȋ�<��{3�N�t�!��Y1�[s�g綱KI�*��|�9����l
Æ�)�qg(b�dTޮ�ͺ=�P��+끚Y�q�;;�L���_G��!�L���� F�5�5����\��)�i��<֫�pK����*Gfk;r��pn���B�A���D̨��5G�3I�d	�&�cj��/�d����`��޿�2ǟć�ɪ�&����G�n�z����)J�	~\��ްRE����(��D�<eU�z3��f�f*umC�C�����QC\H�k����V���VR���$�p�P�gxo��۔����6��_�Sx/��M�o�Q��@ �xr;����:�'?�8�"�<|�=�����+��?�� ���툸L���`r����o��������
���E/x��bN���$d�<dr��}ƳHY,��c ����� ��S��I��%y��*��;¶rq�Ƽ�����dAx�(�W~�B�¦����NAC{5p�3�z�G��*���n����_�\��{`���R<�,���R)_�fC��y�'�$rH+Ï�h��g�U�y�Uނ�x�OV�� ��jjjG�y^�q+<«R��D�j獀+�[B�����G�m���N�t��;?]_y��%�<�k���&-�iy:��3��~���0�J`#����N����"��I�mW>��NA+o�U���Oڱ����ƞ�I>QT�I�%:���j^Lg<��2)��b9��8i[�F�gSM^�v�?1���2�ځ$��O���k�{C"���+������I���X�?���E0�'?�I�<�q�:��I�˼W�C�CgtM�-�l�
r�CC���F����+Ho&��f���m1wLNE������7J�Ϗw���Lh]�n�ؼ.٦�Q q7q�~�)�Ԕ�i���o7��Ͻ�5�@
�ঽ>���1u񁩻���V=F�:n%��*�]��}Lپ�2�o+�����m�e�}����~ �Rr����|��B)��ë=F�����:%��7�������[v+�sl*`{��zH
%y>3t������%g���o���t��-FEUߥ>�'X<1|���TM_�Fp|n�,H�ӼW�c9[�9�H���k�;��tr�X�Ʃ0(x,ry0���"��{�h��U�}�cO2BQ��\+#q%���z<j������Tk>R��|�0�o:�9��m�y���&�����#�ܩُ�^7� 9��k\1j>�#I�d�s�����cB���3:�ekT��y�)+e���D&	�T���=���Ec�8_CPS�*��	�����Yw��q%L�'͢Am�F�(eT�� �v�i�a�'����#�$�؍��ErS<��ub�મ�Xo��Q۷��{JR�ϤR	�#ܞ;?C��r�WF�-X5�FS��{��W75�4x�m�;�
��*�ԟl7��Zu����\ӯ+�}V��D(s�e'֞��3�}��5E�|�A�ε&�&����6q�}�p��K1�W�"�E�$I�M-�֋��F�U��� \�|F�A��+�8�9>zY7�yO���7u��Wb�ݼ�K�i-`��t��T�Y��Ͻ3w��L�H���6��6�-�)-�9Q%��"����ֺ,2�a�d��(��7��| x���P Z̚���3p�n��^�����x��iəCi��_䭺,��g�l�S��si�ɚ�yQ�0|%�J��H�:ƕ�^<?ڜI���d�Bd���8VՁ�������k+�o�Yb�Ȯ��[ ]�Ჩ̴����������k�6ϜE��i=���S*q���r���@�>�?dyg�[�<Q%["�����H^Tm��؋`+��LV����,2n�n��
~�[D2�cl<�|�F�2������&I=����D��jx}?˨�%S�f	�*L���l3{�P�j['MA�ǐ�I�c9S>-i�����z	��{��\Z���H�;���������L{�2�1\QC��͞�DۂG�|Zbl�UsNwZ�����~P�}L#�I�NƗ�q'.n��Q�Y�L��mh}�s�ΙZ\�b����'Bt�<Zp�'�8n�!_�4��&��ը��/�k�☛k��v�yk̐/0es��Q�m���s�.��H��dt�������t�O������m���T��r����)U�s�&��]q	(��l���E/yw�'r�K��Ԏ|���>�����v��#$���Q�?�m�[�(�%�����@�գ��0��ا@je�{�NPờ������ѳ�s�X|v����)�9o����0%���{w�+�4W��1�Ӹ
/WIa�7h'^ok��8Ǹ�iXݔ=�N�QEٛ� ���?����i�����Eq�����,�z�к)��
�ȑ�!�hH��<�p�������_�B�D��b0��������2�%G48}#OP�yj��_|"J��:*��a��f�Wl��)[�<�i谴�芎��cn'*�>�F�6�t\1Of)R0�mb`���T�M����?���|�fs*�`b:�T�w�)��/Us�˨gǣ����:��1�ev��h�f�9��I򤺦W�#���@ P~2���|^�<�|��W�K��^�W~�5�yk���t�9ͪ��j���i+(-g�G��F���K"��t�߆�����sk��s�v�"�&�~!m��|���M+��%"�D�a^V+���:�S�L�&��=A�)�.��Ƒ����a.��*�sy�f[�o+q�z|���#�\\O��p�ґr`���f��O,�!�ӿ��5J��㗬u�i��H=9)ܟi��Z���"���
��0���s79�,X����K���{pF��f?�FE���TR�y�Z�X�!��h;A���G�mb�;��ϙc.���8��s�A �'�Һv@v*������Q���ݳG�<7n�R>�S��P�\[Yէ:��w�=�#y��R'��p۸�Q�2�Jj�Gu�*h�T�a@)�%b��*���E۶�^d�!���sy'���,U!5*���&���ѶV�W�զ9�$�P����Jk��n^#�o�/�́��G뱑���0R�p�,�l�(�w������0�B�lR�K�E� �]�RU�,��Cu%����Lo�����+��q���-U����Q�G�����^iJ��Q�c��!�7��b�:��}ĉ�ɯ��=�+	4J�Y"I �z�J�XP�\�N	}p8�0Z?A�O��ܬ�.�z88)�u���`�ZL�\gS^�:b|��h�&@oH��V�Z�	+=��id.OC�x~�{T�1���Y�`���J;��<���x���u��sDa�h��x����}X�3hlb��>��}g�W#[��m���h���z�"13ri[�b��-��J0FqnV�q _��˾h"b�`&@ȖF�X�Lo�G	���(����������ߺ��x'�PuF[�@��!����-��因�*����"R�lU���<ot� A;�
=������������1Sё�b��q��[�l۹�.�����"~i't�i#���#��}����ᛈ.��A��|�"��k�L�/]C{ɭLq_p>��Tw��zv��j�R����?��}�U�?�>Q?O� N#�.�:����'-+I%8�� �h����1Tc�=�b��uZօؖT9v>��	�F^���'F�P�����~Y,�VE��fr�������B�;1��o��r�?��(��գ��.��AV�ˬ���ⅆ��6��7�`�秋"c����C�%|�g�{�-"�,%�{&m\�iE���>�6Iyv�j���~U��V�rҴw����-������d���=�vRԧƤ��"hٺ�qߦ���_1d�����IB�w{�ݎ�T��^|CI|UW�i��ߧ��e��OT�ёX�O?�Җ/eX㤅o��wR~��6^�X|�Y����E&"���i8�^"����{��h���w�i��g�q��<��V�����X��i�q`���4,�����mɳ'_��L���`Z� �`�QN-.]'D�M�@�A�CT����YF���Ȓ���g����Cot5`��D�)�Y����-�7�}Va�Z�ɔ�_�؎�����8����M��!:R&x��_|],#��+q�����+Ј}�8և�Ι�:��[��~}�o����ݻ'�7&��L8Ols��wfX�Y�����/8�D��_��e��l�-���_����;6-Ļ�/�r�S�<�#������|����u>}���X�l���XD~�h�m���
\��3�H��a��^&B@Jy:c�x:�i}n�xqQ<� OR�%o�wg���eu��W���ʓR�bX2Q�g`�	��-=�(~n&C`{-�hK
_ 7�4�����t
��ָ�\��U��R�F_uG��*lՂa.�n�����[�H��.�n�#�o^~'�v�y ��^C��t���H���pt�V���j/��8�l���\��NR��{V�r�x��uM�*&�q+��E��HqXisq��s�J��X���P
N;�t�=�Y5��_Q7�Ȣ��Θ�|,5��%6#���C��J��$'�^��*��0ԃ0]7����&��`lof��RP��%.�q+��*��U^&��S�>�K{|���TH�����٨.*�ߦT^��������k9���R�:UH\?7�BՁ��c�{i��/���l��n0�����}+aKC������b}�%w�����+���,�oѨ/oeg����R�C��L���}�R��b�g�-��g����/�p�R݉�z�'���o\�B�dK%�,-��.yz���R��Q�Q�1�]�HnN ��G8��(-�=��o�zm`��()���[�������~On�ġrG��_.6�S�^���iN�+������5�3؅����`����8����K{b�b��%O�|hC�K�F���y��k�t�甬�Znq0l[<��k�˘1]�}�?�,�_�s?
pe�f����%�<ӚZy�f�g����[���蘰���<Ƿ�]N*�d{f�kp�d*ۯ5�G��a�?J���|P���G�v�����'�T��������PV�J5�'���U��=��i���X��2��É�Qh>��5�!Al?�� ��0�|�� w\�%X�[�z(�Q��Y�M$a D��l�����(	jN|��M0�_�b
�V���a]��w,�U��\V��Qa���vl����ds �4!�&���N
,�g'�p��e新Q�]�Q@�Q~K����	O�`LZ�~��s��U�H�i�[�B���$� =�O-�M�p����7�p�Z+�=a7s�"�����6*"�2�ݷ%+P��R�
��������k�*����5q�IW�(�z�5�"Y�x�/6�8c9�#�<Ȱ=��# }����'�ǌ�CF�Z���I��"�k�g�L�̮ �X)���e�����Tn@�!�C//땼�f�;��CS�US;��i�l�K}��}�t���guayb]�/�Í�gqq$1�U�59�����G	P�ڼ���5U�ͤ�yV��g]�ac\z/��h�����19��~H�� �J](�m�HQj�\+�����ߓ�������h�Н,3D{��_��� ��)F��S%������P1���I�e��Hj���<K��:ϡ��E[�a��7>���E����v���
��LP�/�3�g��&3F��)Y}���h;΅��s�铮7)�
���#��䚬�˲5����r����]d��uH`��vn8��{e���}k=G������Ok��ɿ'��] bI�?��>G�{9�=��^K��	�zD�:��h �O/+h��DP����[\����I�֤�S�e!9�_y�/D���R�}Xs�V�' L����.�_/�8�X��LY����#�7P���A?��|%��;Z�D�N1e��e�T��Hy�J��rcT� |���Uda�^L2Y�cp�����k���o��V����6E��kЈ^���xTv[��u6S�<�H��!}e�"�ɘ1[�f�{B΋����^zvրT���ڏ� @F��ͲmS}�x�� �	����Rh͛�X�m��p
���!��q��_�ώ���%�2"K��XL�U�(Ļ�L�=���U��[��b�r�L��Y��]�G7�ߣ����3')S���]�Ϯe���?M��M,ͥ6���v����L�2�x��{��x��B���f*
���(x;0�l��#h��ζ��I
3X�����
� Է#�7�uc��mf���� !����� ��T�}RDU:.�����m�-��t�?;�4�#���7�� �7�xW�G�f.D�ց�K��.V�����o����U)5/����Z5�;$7XE���ٷں}�-�\���N���rl;���s�� �;b�gܒ�����`��Q�����.�%�7�o��!��?������r}u�(S���?MZ�&��AHCf�.7e;zc����Qc�p%���)�nĕLvC� ���\�*�o�_~?,y���n=�&e����5�=�>Y =vG��9W�fh>����$r�ھ�z��I��Z���v��F�Cg4j��h~���Aݴ�No+\�S/_Ư���`�?|C����!��XL�#��H+%�%c���M+��D&�r�ǋ���"+�WFb�5o��s��u�JJ�KG�7f��к��~�;��}W�I��Y����P=	�2�w�o�$y<|k�+�;�4�2ݤ�2랬����e�Ro���lIJͼ�D�7&\�l�`�������> 
ӣ��ձ�8�?;o����h�{U�=�Y�m��U�F�JRFY��a�Tk����y@�@��U�1��N{H�mq��-�1O����=w$J@냔M�j�W�/KS-��.�M6�u3�&:؀��� ��n�N*tc.!e�4|e@���JH�t�twH�4H7H7K�t��t�tw7(KwK�ҝ�����w�`��9�Sg�u�˼����s���}��)��W~����|ȱ�|�#	W�8�2%�;��O1@�!̱Ӹ���f~�:��Lx����)�!�N�u�nSMY &����C\$,B�D�ˀ}���0�l&�>&���W�
�6�h�v�j`Ye�cf�w�"�-BwT�X��!����Y�*mX�R�/�����,	���h�L��g�oC�<��!;q��1r�w��=��ʷ� FS��2j��VC?����p:�od�p�+!Գ�aXA���])�A��&�͡���qH>��x�NŸg|��8u̐�.lB��p]�!�?}�~1e[�Jض�{W DQ&U�J?�?ݝUWX��߯�n��ڭ�Us���ДIz�>���$��%�<ƾq0�Cv]!���$^����EX���TC��&l:&v0^��!p��\�'���w�ya���Ir)\�:�5�  A��[:\̘��8n�3�D~�$o�"�����ϳ�ݱ�j�ǈc�z�i�1�r��{�r:�/����C
�;ċߙ喦����!%~�&U=I�FZ�z���:ZY�*�К�x(�Ho���0˾C�#&�������L�xf�8C�O��?���s�K~���������zu���Ҋ^�4��X9k��v뺟릈!=*�/	�����;���pV�%wh/���d���V��c��"�n__���
.s���O�,��7�4��H?`!+�C1=G�*\j�|�#,��ꘫ���=���{^�im�[��r�m=��2���dj+h�Z���I�i����e�@j6�s��6��p8����H��}93����5�1NTݢ�Sst',�զ�	�
M���� @1e6Gy���F��Jl�ϒZ��+�11dΈ�#~=�J�u�ݯ���܈ki��V�>�~Yw�ņ�-E2�$5˩��Í�1���L��nN��T��8��u*d;�$j�bP;KTM�<��^E=��g��X�oO.��?����t#dȕ��LMULN�5��:��������2��\/!��ө��_3�-��TW���~����&�rmE@c�|#3���P��!IA���"
�b��8$���˫��m�#G�� d���.|U��`�Z6�}!�!�Ib<W+[�@Fw����jr˪�T�
 ���P��:�M���p��u��@���)G[NW�΢|���mtxC�O]��Gխh'sHט�eR�
5�[9��쀶5�������#6��۫:ר$���1�ON ��� �K�:�� ���ZB��զ�F��i��������£rs`s�z�J�M>��X�Y>؀�Oc��ll��
��jѓ�|��M<j��5f��	����5N�����=,�{�����?И,:����_�a2n�h̪���A}6;=�
*�1����f�p����2����y�d㔄^���<��I���ɬZ��5�� G�#���G�;��Q��X��k�<ie�`Z�������Ц5j��"_�6<�xe'��UC�Q}�U1O�૜zg`�D��ʐ���!n�Y�x��Tq5�t&��<5�l��!z4�8Ȇt��]��S���o�(�Q�D�T�y����Y�h/���7PD  eS&^���d���[�X=W�o�����3/^���U4fr����u��w�Ҧ �s
Ѓ�U�0�����=zy1c�ʓ(�MX/q��H%Q�9b)��dF�DI=�.���y� @��b9e�' ���'��|l颬�8o�p,7�g�	��]b͊��g�jY'0,  ���~��%XϏ�Ō��+�Z�zW;�C<;W5���3�-��3��C;N@P�r����r��*x��X�5Q1l��1�����,D#��Cd2�d`�SnLDEE�73Y/�Ӵ;d�Q>{�M�\��l�,�쵕�p�h�p  �)���$p�t�<}��^�ѫ�D%�qs�/��2��WQ�����$�4����K���a��	]����x�{V*ܓA�՞V�~`h���B}Sk���F��d�|?���(�����b���wv�����G~���% c�`�~�����O �i�4O@���s�?M�,D�Sޏ��d�p��H9ь���JگJ��\е�{�������j��l8۷J�+�+�i!3����K�0u������;z?r�����y�
��(�o�>�!��B�[$k,R�>TE��;�4`X�heεr}2v|�j�	�����܋#H�%u�/��+s�٘Τr����d��Q��>N��l$�}BZvٲ�Q��S!\98%�\�g��p�I�C�O��l��!�t"�\�**��K|��֟Sr}�k�JU{53e["��xb�sC�Y>H��վ�\g���鸉yXT�da��B`>=+� �ҫ[�lq��F�A��%��/NVj+H�9���$�[�='��HզpM7���l#WS��@$�w �w��nrݑ�>�WͽU�#dqĩ^�۱=�5��`�u8�gy"|�1 �����Iֵ��JXm8�gV2��x���{S�zhI͝Tme`Cm �8���"�=�}��+�֤`b�k�:�m(��k=O�=�<�I�N1��X��"֦k�wQo&��{�����%Mg�tOg�L�vu/����	�]�P�:FY97Gx�x^@�Pa�V�Q9�&��kw��R�}�ޤ���V���\8U1����?�t���yn�����?��+�jS���W�..���Dy�e �E���V:	&+�O�k�-m���]�&H:�Z� #�n�eE�iNnF�u�r]"��.���p�Ig���rqE�3W�D˞Mە)�@9$:" 5��BA��,���
��ks1���ɪ? �Ҩ�$�D�}�,q�vW�6�O��ȹJ�8�q�; �������G�+kNx���4X�۱r���6w3�.�X���Μ��10J��Ic����Ma�(�e��$8,2uM�~�a*�D��+���  �|k�na f0���P�ZRA��������<��F5��|�p��~���[T[y̍0R������uW��r�}}(���85N��!�VHf��
>6uҠ�E�jW:Y������vcn��L\���JfZ����dSA�uP��r�?d�AJ�Jc߿o�%=X;��=L�rj� ymY�?zvO�T�y�$h�B��sUF�7��!�^��~�/D��`���5�/�N�H\o�S�`�  ~�nV
)���ΰ���m�b���5�lK6��q�;\���?��!��UWz!(���̄����\���;?�:TW�jʾ��`S�3YuJb[��2<i *�x�r+M�|����r5��[�i�����I���z�c�"��yQ�����jS�F����t�Y�pY"k�!���V����G'4���=3T +�k�K��i@�)Iԑ"4`V^9�R�Uy���e�Ңs0���.��s+���s2��!2W���[_f�PFg��)��ՏM�/O��yW�UE��6*U�6�����:1 �d�L�y�gJWB���Q~k"���-7��͵]��a��[�E�N���cH>��/�����Y���D�(��E��B$Y�rnL�~���oZ�"�ň^��=e���x�� �Ux0���w5�Lu��~�;*A��e$l͈ni��&B^Әh����_��Q7}���<7^,�U����C
��.�34�κ��]ٔ�deJ����f+�*F۝�l��O��G��W8�����vԭ�Z� ���'�/Dc���O�����8��d�f�~-[w�m�s��;���eQl3y�b�.���٨,�3�#�71W�m6B�c���6��h�rz
����6�����ۆ0~�ɚJ
��v�a�:f���B�ܰޭT/�[Y�8a��עU����p�/��>� ϛU�K�:_�īZ�C8��hL=)Ơ3�X?Kz"�
;�C�M9�S"4���0���iB8F�.�ҽ&}&�u̝��\ߢkP����|��k��@��МP���^V�h�]9(C���֌����4�I�am���-:�����]�j���sIrsS���D���r���n�� �b�� �+��\��O)�[���UАm�4�R(�	PcqhUsM3�����r�F�t�~�͓:`�`E؅�}�!�vn�G�qpa��BJ0?zpu|L�J��`h�'�x�C�� �ʫ�9_�
|�I�~m.�����=�:}�%�����C�3�A󡇄�#Nq�h,!�_��C��TY8��v���E�*L���;GSV\r���;�hS:��Hxn��-P��A�S������g���|�0��â۽�z�g��g&��? n���*j�)���q�V<�Fԟ�8U C���L\Z�r���V���22�4���m�,���{�_gLl	r������8�k����t,)�1`�P!�-~&��<_�~�8!7��me��d�يh�2���%�mc��w��K�HF.+�����ZL�s���▇(��㞌� �m�b� �ӌ�>�b�d��Z�_���h��d�7��Z�yl�;������n)����r��7��"ʏa�NQ����e�q/;�v�`n�wYr�[��YXM�)u����f���������;����BH�Ϻ�?(��,z�:�x5ECe��V�.%Hs�6��%@��a��V�0)��Ɵ�y5�6�ϲ������zIR2��*1���o�˜o��`�O��� VJ�	mS��㮏��H��4ޞ�4����OUh�]cu�=9�8��@�٦��2��Ƹy���l�9�#̳�c�����yL�-iN�����*�HǵqL|�Y��r�t��6$-SS�i�f��D	���{��	N/��	�t�h�?2-���D�7�����%V�=�zT��u�I��K]$��ż���&I5�aI��b$>p��G\��6ta��!��u�z/4 Ky�Q��D*����J=��]�&|X��"h��x����.�?Z�2�N��t��$��B���&�?;[-Q�SQ�".G�4F�1T��R[���i�-]�A:����R��Q ~DD�0*��d+Oy}L�����#�vD��=j�m�W�H��𬯨<�u�,'��M��BJgޚUSr�#���?��Н�/CO!4(�boa���E�k�m&��$j!F�S0=w��e)�Mƶ��||@�S��&�,�����3�[���P�`�M1����;��u�׊ ?��d=�$�N�	�v��5��]�U��]DdvtKB��?	Mq*�ƌ蚾�	 y��L��D9ܧ��!K	�,jK>����-�:�/+#�&�&����O2D�>:�$���7]ߎʖ�N1����0��7���<��9�/Q'�.�|�Ñq������z&�v��ۜ����| �X�'��y�3U��<�r������`|���8����#��5B�c*�6:<̕� ��a���~��Z-T��$�v.��޾"d��t�q����`�����r�Ӂ�h�e�/�@���0c�_���J���C|�;
G�t��ab�(ێ7������a��L�R����xY����ܼ�QΞ$=Ħ��Ε����[�ݴ�g�n�ʵ<&<L����{��SX�.6�Y�i�HHm��;>W?�Jm�u��l�k�=��z`J}�A���r���I��ϛ"�����6^.FF���"��\�'	�� b�Ub>����\��\�UQatՑ����e�WP��9._��cJ��~�>\�|D��7�~��Ј�'����}����l!,��jnEOGE��&v�f���s�@f<��	a��+r"�Q�&�(*�U��D���䃅
QF!_qs'��~�[�O��Q��i��:i�Y��3a��h���f��Z��݀��%����I�d�i��ʊ.����!���J�0�e��{Ӥ�p~T \��e��_>�u>���G>�N��W�d�m���d5���@2��eVy�v���K�v�����(�Mxf�J��8���A��[h6$as�䠵d�0��IUչRl_].Y�V ��;�]�] {�o�6+`���Ԩ!N����<�)66�MI�nV��aᏺGV�}ɴ��TM7V<����3"�?�jߌg"�@���.�i�|�]�]�>T����=��5��4���7XPc2�9��ڒw�EPa�G��5���Z�ݓ�3V<²e^�4���9�eo�K]1�����݅ޞ���}',�|�7$�=���uu��~q{�d���������	#9\������8��׃~���#/蚻��`[o��m� �e`K{�#�g1��J!C�Z�Y����g��tg+ ���`�$
��� �lC����8�v���N&I���ugZu:�P�l]Jx���×���|#�4��h���u3����t��!�AP�D˹ut���#<�\�Ʈ(����0���������M(M�B�i���j�H9�K�ݣ�r´���˔[
�2�O��#�D��L۱aqs6ߔ��^?�yα� ��OEÂ���r�?q��إ�W�&7��g�'��Z���.�W]����q�\#>��x�[�|SB��uS~6��Fk#�=,���ƪ�"`��{�x�̔�𥋋/s�=!ꗹ�Jh1�o�؍0��������r��9�PN�7�2L�����}hS�=�R]��C�Y�����Z���>&a�T�C���f�qm�H�5�R��ň�A�x0v�#K"��)A)%��-<n��'$u	�9�s(��F���y�zD9993���]���Xֻ�dj�2���ˎ���s�7t������]!�=r�/��韐b�#3 ����C��`bm�s \�5q�.�5�'��'���=�u�xc�u�ŗ�Yb�� ��Ѭ�82|@�OBJ�y��8>�r
@O��[(��n(���t�;�������V�ǘ8ʦ=y��<�U���z�_�����(��kTC�+��"��l��-z������<j��Z��C��M��1���Zq��h��,<�Q6������x�����`j��`��Ҫl@.�G�����ˈ�}vJj� ��I��඙�4!�/�}\�c���.H�5�+�m�ىD��Y9q�0�όrڲ�����GU<?�a4n�l�&fs�ҡs*kҚ����w����g�)'����u5�@ɒ�Ю�9�'.���@�fb٤n�3��d�q˕ψ�0��o9s(H$�������)�n�dO�ɍ�v6~A�wJ+Oq�� ��0��2�������&4)�w�ìGX�H���ۮ�	�@H���V�-��B���c*�������?�g���wY-���i�OXb�6�8'��a��� cY��=~��e�󚹒�\<{���Mt?�v�\`��U�����Np,߱*]��lb`���4�*�Yy�d�� Ëf���O����Y��p�%-.C���Q,����JW�-U�Z�Df�zg�w�d3"aӒ�S{�4�95������U��t�����Ͻ!wZ�~B�#q&.F���,��J�����@��Kn_��K�yj���~ۖ��\A�W��zJk�*U���zY�K}�z ��a!�u[P�%+�
2�"����5�2�cd![�g2�Jw�!��㝿���C��b��|��2c�0l��EbnW�����}�<*�#e�����®W&���x/�9:sخ鳕" ����!����K�>ʜ����q�q��e���ծ��c{����f���u^2��`�8�a�c3���׆U�"c�hϔ��p�W�Q��M!�-�N��F����tM��!�`6�!�𜧣.��5F���R��*�߳+���{�X���m��8_�N��Ʌ�(ZVl.�/%�ǻ����4;�2����mh#�?�=��:�����|ln����gE�E lo7E�Kn� ff����r�/�����x�g؞6�W}ѧnk������oM�HmO3��O<�����il/=[���Yj�g"���bj�I�exf�]��_,�"��I�rֱ���f�r=�0�m��B�<<.�G��Hi	�v���k_�v���d�ܼ����T�U�U7���q�v���8�&+�bc1�;;�w���FCz��n����y����ll-9n�bMkIf�A+��=}=|�b�)(�C
1Qd.�~]�\��9��W�6)���P���%��&.o�z��G>�&�<�	"��
���,�?�S���5�7`�6�������-��|O$���� Nωj�Z|�'�z��-� I��2Zs1�����ܐ�=�o����%�n�aP�]d	B��� l��S
p�1H���ks�#��J]��Ϣ��bm���ӝx<�a0,T�@8�?#9=��ys�}R<�!,r��6����l-���p���?�Q�T␦�����G~z��HI\ߴ	Zs醀%t�~}�\)��"h�R3���6���l~�}�ބN���G+&��r}ε�þ�_�L���F�>��2��'��(�簶�8�Ρ�5�#ƫ��v����¯$��c��K��N���A8FQ`�e��٘��5Z�G�T|��Z;( ��j������ܱ��[�=�~@����٦Jõ�ġi�krv�Ru����I�S�q�@;Ih�J���ECl�K������.�e�LTz�t��K��ö�!���F�*��U%=§�.)@qpyb�G5}0ƕ��'�2��K.�Fr����d.Gط��Q��`o�����r��l6tS�qє���aV�?yH!L`�}�����l�d�|Q~2�i��׮�'V�_���8��<,p�i�y�n�u���ڦ-��[Lک�e�;nM��j��L���H/�E.^���oX����� F�x���Z��/�듢=����.ć�@Y��7���so�1W�H��(�D��><;qHc�/{�ɻ�q���u�>����������<�x�m�W���§ѯ����:b;��+tv��gxy%�}��3h�9q��yOe��[��~%���c�VF ���%����7���]�<�N�h�e ���5N�}�+�}�6�30Q��}��l�m��6�IF ��wk�׶��y�_�,�_��ݣ�ӈ*m�ɷ������#�0=o<9	i�VcjI�w���4?�@�m��D�,z:b�f�WP]�����%�!�[�2Ǽ44*X��!����itc��;v)�I�kʝc��)��f�Z-���w�w*SV(�ݴO�w�ɏ�G��i�bceڏ����C�z����Qi%K�p�.���N�/��!����:j��*s;���S���%�����\���L��$(��1�]@��f������K�p ^^���y��Rb��d�d%���Y5���?��a!?	E9	P(�d���%P�;g�2���e�U�sO;��դ��ǋ��ǻ��q�0�2m����w>*#�<�~ʨ�I��U�8���UiB�x<[�4�@���c��x�Z��=�܎��UƳ������n��`�� �s��d&�Tȿ8��J\rѨ|�;#(�k����∩�$Y��y�e��=���L����f�] 1UÏ���=&ˠ+<�'dm��}�P�@��<���^����0��r��"���&AA�ʵ��.ݯ�����(27��r�uƟ2�zm�����r{n�+f�S�������.3�l�f�Q麁��}��;#��AO%_q>��ʱ-42�V3�w�}<v,��J)��������.�!M=����"|���RƫC�ک�B��c`¶ɣ�&�'�V��ח�����
��bA�_L�?���]�`,΍��tM�����>��I�H�7���x�]l�˗c<�������5��U��e�.!��!��J��T�m��w"�;�a$��I(����&0u�`!��#��Qy�k��(+F��E5�l�Mn
r��Q�yX���(����J0GRm�
�s��g�[�t�b�ik�@"m�O*��V��" M�8���G����j�����ދ����Cw��Y�""���78p�T�0�{��J�?���du,EjO��ё���p�B���z!�J��WlJ�G�z}w��?��-�9��+2��\]~�xY����>T�:�i�)��3g0�ieVmTL��6���U��J���͋@L"&�����R�{�&5��8�	��I�� �p�>'�I;�6����~A*f��Z��]D�gk蛰e�Bp��&�^�Ե��P<×�˒]O>R����!
���e /��"�]��v�Lў�ڜ���̐����pe
�E���%���u���eZz,�\��w"������u��,��{;Z�s|�Ņ���/б���$��$9�s�a�����O9�?+Vot{��+��%y�!I//6p '���>�jя���m6�(ю,ŕ3��I0/w�=6FS[�b�p�|)ۥ��5�D��A���2sQ)G��*Z⿷/�^A��jd���ǝ�KSG�Ŗ�
ĻN �������4����,͒ݝ�s�N�;>>^Z�3]�<�9 �ٔ�̧5B5 L��˖����>�L6R!v)� ��`�/�·����xJ��a%��0I n2%����Ѣ%���_���g�6�F�o^��Lo�Dp*$�R��NDU�*�$����<^W�(/���&Q*���y���{E0L��>3*S�r_	(Lߦ5����
���[dǬ�?ظ=�<�}��x��#=8Y�\^�^j�i�$��i����bg� �^8\��+���R;�֫2�>	�Zh�]�~�O�9$F$��C���ex<>�>t���ɚ���^�����ܤ3�K�q�&9��|$!a��v�/`>:��-Z��w�&@�Su�
âs�B�jɋWg���5�h��/���\,��}3fT,�3��U�H�f�O�K�E�Z[�3��n�]c�2}����˻���a�Qk��vN�2	���TK.�]c��(%Ɵ}׋YGTq���{�y}�b�΂=	�Ig3��Q[�? �mR4.���Mt�M�=	���C�o�n4/K9l��z��*��ҝ�L����35�����|�5a����n�E*�_��Z�v���]&󐓓����m%T����n�<�D�w�gY�z+�D��M����,w�������N���s5@��v-q9�l���.�ܖG��;o�B��L���*�������7�>>�5:$je�=���� s,����E!��>5J���.�����Q\�Ű�Pq����m�)��������R�(�э����Y�ܸ��N�����2�b�Oi� R�ڍ�R�����"�����	Ȍ����`�P�.�:�|eRi�0��q�ۆju,؇x���{x�eS?Jb�w��f���5���+`z��	5�[��B��N�m��K�B*����VO~��~M����G;e~����������	"2a��#~�.�u���i:�b%2�v�y\U�=��j�(����_ʅ E�@g�~����8�vem�,*|�(��C���H�$f���ol��f5ϟ9�;&?f�6�#�H����,�;��l�]��xw�m�1���!��:.b���e	�l��*#:����5�Y#��l������� Ph������9
�[��y�%���4��|q����ݥܖ~淤��x��X���$rf_#��H��T*V�G��+rM��E�b�Ҙ0ݦ
�h7�����ɿ��A�f��1��6P�1_��|� ���mg'8�nC��)�j� O�C���V0���ٕ����]�"VQfӹ�Ӷ���d���Va��=B�����ge����%쎨?��N��� O$��kH�i��Ӛ
�:�էG����F~�֧�Ҕ��Ƭ.�qV��g7�_�q�%�}3����g����	��t�Wj�J��lR�������g�;�|/F��'�hq�>Ҧ��bc�gK/3�8Ӥ�h�T!<O���o����e�{�rF#)m%i�s�&~R���d��^�yjH���e�	*\��	R��������s�GG�Rs�,�����	�hMQ�Ƣ��d*�9Lw��vON��<�b_��м��T�m�;��:�A�ӫ��l�)i�m��x�|���U��CUa�T-�[H�3�WD����z/i���ұ���`�G/'�������1cZP&D���6]�6��θ����� �E����Ӻ�;>���@�>�����8Cۥ�&N��.�Ͷ)������lcv�h��z�:0p`E(��V$�Y������a?L��Y��:��>A��Y��oء�M�\��|�o��;�^�>J&Y��F�}�b���aV�������k������}@��]�4��fld��J"�k�9��)�Zz,0��4�KU;T'�%c�^�G�y>Nfdi[������ӢԲ%����li��_'�pҤ� ���v�ϋ��
8f�U@���Y:��"1�������ޏ��pr����\��=eno���0�1~C��81XUX4\1� �{�H���]f�� �g�PXp1��H��.k�t�1�����OO���gH��9�G�c���-]��];�qg?����3SCnW1<o�ħńc٭\W�~Gz.���0�%K�ث%*�)�P���t����b�s~��.s-�M�����ޅ;�kG3]ot�"S����Yj�s؄��%�P^�y�7p6�������<��ڌ�0c��ol˭���zj�m�$U��U�T�/7㘰��5K� Ca:�A���K@�����m�Iv��-�텓�"5Lg�V/A���̟z��#<�
��TXc�\3hid�C�t/��i&���Wn�
funÈ1!�;�frk�����R,�tq������%l�,����I�f����N��=C�'���%N��*�@�1*�����Z�Z�ಊ��t��Yc�C��:ר���.�	U�Ix)��,��2k:{�O�+
B��:	�ъ;��b!/=3q��L��a��y�FUu��{ !�ok�v��S��j���,�;��.��;]-4Ϡ��Y��b�h�F~�mԬ�!Q�D�?��P��)�SXц�z���Uot�"�����L.�]�P��/	ᅝZh�Y�Led(�X�?9u�,�/����
������bfa9]`q���%F9�(?o�T` ����4�L�V�Ԧ��o}Oo(�Է#84.-k>X���N�۶�Ny|�4n֝�c�>s7@xi�����Gn���N=��}�q��һ�� 7S��=t?�'�$u��~�d�a�E��7V�X`�e��r�\QA���o�H�:Fb�̌���lVv���8����R��z�@keX;|��'��+K�,Tbb����'Qݫf���cP_0��C<ox�i���:�`�Z2��Ѕ\Q�S[k�4ڞ���p^�?��f�oծ�LI+��dHP�l�%_����H*qV�IR�mC��7��K:s2�}ۉ��R�%�è��H�K8�e�)_ ����<񘧷��O��@oX�"&R&]�<Ggg��i��B�%Kq����&��R���7���(
Gni?�T�G�񭁗!4]�}e�h+?�-l!�����p��i`h8sw�qx{�rj��#O�`j��k���h�3�1��-���c�^����)��Mo��UJ[�1�#2Z��s�bQY���ۇ�xw�"���>_}�խq������V������ �c`(����Un*�����rSTC�8e�D�$)׊"'_�kD,�7�B�/����i-ZҲ����`��}_��_xV�>P�Ѹ\��)�+��[dR���}���<Fk'k}T�����N�sf���{�		F	�R|�d�qUq���0�"��^V,��iٯVV~�.ƴ�t���t�U���eEP>����a	)��[�R�
�vٛ1�ǉ:�E�h+/wn�!�fAqY��jU��UfC(����׎���t$��X�X>fk�����C��}���VD�Գ����Fzg�	lZ�4||�&���1��w������(�ë4.%?��V};� ��ѡUu��^c��q�@a���	Ż��%��?��v�B;m�ҳ`���0�들X/�b�� ���	�w#(EV7�����Q���W�+�A_�nT)O�揃÷�����C\�w�����I�ŋ�*����a����ܨj\y�TyL��oeO=��S8�T���P��BCz��{&�p
)j���"���o�Z�Ʒ���t	�,�N<m�8����ŵ�O[W˴9E�U}M���+]��k�5���38";?Xn?AU�EG�ǟ# �C�*ܦT��$�,2��mE/�h�aL���6 g^��ww���A/Ш�3t�K*q�xi�}fIC�0�[��m�V^�tM�1sxm�y��cg�DG/����*z�����2���hr�,S�4��/���u�A��˪JG=�;Jg��ߞ�6�fWi�l5���W�җ;G���>��;���?Jw
rIf�F ��:��y��Ԟ<ձ��B{��u��ב�9����\���ϰ�V�sT=8����QP���$_t6�+�B�ͺ���5I ���M����5գ�×ǋ_"O�����x��Hw��и]�v7J���;�|a��k��08�/�y5G�[B5�+R��L�.+V�*���F����ťy�/��Z�䭘)��gc��y\��d��T�.�K�Y�:ep������~h��>�|n �jj1(�Ii�ww��j꬗�>*ǣ*��^��!�YQ��7}3���R]�-��8��
�X��4�3��y�����%�|T[�}�<����l�oUS����o�F��8%�d�Yͪ�/�L9��OjU��8 zX���U�����P���5���F��5�z�Ϻs>����{sU�I�����YU��%�����K�������O��,�z�{�6�P�c6��6��S�!��F�b�/9LJ8�#L�E~B5��I�&
��]V�6fe�8"9�#j���CRj�0��L��X��-�Gc�\ ũ�]�j����ڝz��r�x��rĴٍ}Mj�n�z�y���m�������D��sM���;�a�
,�_�����x����׾��"���\%��}���yp��_8?v5���L��ro��_��ʾuW�Ɔu4��~��
�Ɨ�}�ڢ��/�2���	���I���6d�[��4�p7�e�8�z�4{.(�blp9�6/�s$H�?�:�u��
E�2
ӷ��S:0�Ӽ�1Z�6��(�]��΁S"��CE�EC�°�!l���;��C���(\1���\����9P��UN=����%=�"�19Zce�[�|�?ƻ$k����k��7�*8_��٩�G:&� F!���h�,h��/ PN3����e�@^Bdﱙ�jϕ�P��$/��Z]WA��/��Q����:-p�`q�h������Tǆf<ESꏷX"κ���2�蝯+�q�W��Ϙ���G�攎��_���?>{/!�Ĕ�c=�5Mk�4�#5c��~uRlV�ߜ7�K�۵���'SW�U8ncI9D[%��k@�+@Қy�����u����h�c�R<c���8���4�e��
=��5#a˃���9��E�n�n=W���h���z�b��ǅ�;4Dꔴ멈i9����Mۈa�5�y!�-�2�jӯD�^q���D�]�b�,�e������A��������0����I¶I�Rپ]Iaœ�Y
��H�j�ԁ��۹c�0a
��#�#l�2bev���Wwyvl&'��F��;w������wG��c{S��yb*�5��;�+˄�.�ug��ĭߥ�4Y��5�z�h��I���B��C'B?�������MJ�s�)�-Ti�¯t���p�ǥ�/z�Q��f�Nh��Q�L�sv�T��8��<\ڨ]6ś�(��g�ּ5&^�w�n��FW�o�N��Rw[�c��fj�o(l@��g��\QOE�B����R�@��3�+A��;�Z[)ũ��*�ʠ�C#, [Cq��5�����Q�A����}f���T���4����n��C�e[}@eR��b���y)O:5h���&7� �=�����PO���1�����:���;�\����=�ۚ�����
x�v���1��o��J�t�`e�� �j��7W7߆b�6j�>�XV�|��O�����Ȇ�+3���;8�
Pm7>�֌����I�����T�l/~_Z�<k{Pd�w�F�iɑs�x���Φ*��G'[�������ߔjr�e�T�ʓe��,����]�K.J�Ի���SާUD�<4#jL,1��~�8Ȟ3"�M�k��&]ވ)4�d�����l��N�t�����2WA@�{������;g������4WX��Xh���Nmz�S�B4�n��"tI�WO{��Y�)$S��eA4ʙ�k��I��;ڳ��C�7	�{~�d&��x�5�C���7�.V�l��k����y�0��6Bn��l@C5���Z��jc���*���Je�[;-�Q%|~�}������jβ(k̭�'�cQhQ�+S1��
R�uSȬ�+l#i�� �Q���*-y�|JM��<��A���B;�dg��.æ��*�O��Ǆu]��cت���>���ʖ��s�3�콱5ו��	V�Z�����,���<�g)֚|2c��dJ�z��dӎ!fL�Qk����k���\㬖��v�:h�_�F�= ����;���>z�ȩ�>�.�<�jx�Bի�G��g��&J���Mc�\�P8ߛ�y����ʛ��G���Ek"6�d����|c7��'�`�	����	Z�-=��1=��{p:Õ��"a�jxR i+�P��V�:�(Zñ<��
�@~�l-��dc�6�<�k�XϞl��+_I'�Ѓ�1�������g��PϚ�E�%fl�h�"V3��}�hF���Mk �Mw�q�T�i��ʭOl�<��-�i�<�G��"/r]�T\�݈8>`����8:N��3�j�\F쬫�
ZT�gy��,���U�#�P$s�Ym0���~G��[a��H΁��y�:��~��>X��}�C����1��#�վ�����l)
q�(ʯ�}�~f?w1kw[��{ٲﻇATi�����:��7��ڿˮ�]}��0�mM���L��������`v������}�H��½�f����u��̦P�a��ұ�"J���ugԤ-f�̆(2!�A�ʿ�H��~+���C�=WX/
^�l�����i<*�V0Ya��������5m>RW���h6�����6��G�*
d`ñ���g[��%���eWǺ:�u���4ֵ�#���"Z�p��'�h�)A����ۧe+�w��-Kt���o�_��(ٞ;~fuͪe���E�1k9����焕�3-n    IEND�B`�PK   ���X���
  a_     jsons/user_defined.json�\�n��~A�-�!f���/k�٠Yǈ]o��X̍6���JT�i�����z(ɑm��tK�H,�<ߙ��}�B%����y���i�sLy1Kq<H�eQ���ь�;˕�/]�_���݋wS����È����2�*]���x���hvt�5{9�Ϲ͝ՆP�$BJbcrD�d��>P�k;�ͼ��Yuq�L�~��{Q-V�g�iżڸ������Z�� ,
N��@N���� ���+���ls��1Q�7)� o
��$5	Z�\s�pw7ݸ���ĵo�������u�O����,/�/>�g���b9���G�ws�xF�
/�}����?Ȁ2��_͊�pU�7�Z��6��eQ��XL�w�Ɍ2j�����F(�/g�\��w�7u>�w�����~��e_����t� ���. ��5�� �@��V���>����/� �@�]@��.���}�j_wٷ�OX��. F{#�Vۉ��"�)�"�7�^3��)�U+��S-X_�x}r�ѩ��`@�"�N�`}%���:V��i֗��]��f�y���:��zSx;D'��7��"�InPO�oyўA�����˺�� Mb� ����C�&�w }wv�H�$��w�f+hRz�;�v4	���5ֱEM:� �'��,M2� �'QhO����=��I��r�$
�y�w����ʻ��?���P�]t�Ay�.u�w}�ۣ�w�w�<;i�"t��yv��E�޹�U�
��;s�PmZ?�7�\���i�m����3��(�iQ��e�����M��S5Z�U��3{��I�L$.hO�"^�D$�2w^'o���{�쁃��灸<Z"��R�Hʭ!j��ؘ=�(C�UNtb��1!
"MO%sx߷� cR���1{�����F{Z&M�F9� ���E�衳0�g�n����^�7��'����^ ?Wף���Ň4*W�&�߁x:���W@��f[T&�7,/�?����a~�Jk�A6�dc���D6�ʛ$�#���-�z����ue�BP�q�Z�D$Éb�s�k4�}�a��9I�V"�1�&仏,>���*<��階[�Mݢ�j�l�M���ijlŧ��D��� �o�7]��T��j��_G��
m�0-�/���XT�+�ͺ韫�֯y]o��_�E�=ߙZ^���f�����?�>��b~t�ϸ�?��闍X�tυ�wᗫE��ET�rqo�����ߚ�|7w����Mջ������U^Ϊ��_�3�&�9rT��ғt������^��(�I.c��-ib�6$�����ޛk�r�����>|�<�����_�}����OoΏ~�ӥ��e^�K�]���;��#���)J
��ҵ
>�dI�'�'T�5Q&p&sƋF��%�	J��7�z� 2��!x� 7� _,b��~l���U�(�Ln�إS�]4 fy�[?�>\�N��������:ښ�)�u�U5����ǣ'��B�-���y9���(�EHO�N��!�^HU/�f.��")�h�m��Y�D]� ��)�`�=l��s�a�7��~�9�����ht��ϧ������(&le��HH��MB^7��1 �J"�҉8�8c�s9 �:�P"�\e�JÛrb�NF��@7غ|��uC	ܔ����mb�f\p	ݲ�Ͱ���b�m�4cc��Q�rU,T11h,\Q�ƳJ�@��/6�,:�&�F��v����Q�I�䣉�7��j���yd��JO��K^���HFZ�6��UTbA�����@k�&�`�RуE7[��~�
+W,F�v�=����c��T]o`y�Վ1D��@�Aup���F"�@I���ZQ11aք�l��I�rHL�XAf��W�,��UJڢU����6C�u
S�)e��jg�+���������W'���.^��x�'��w�S�	��
O+g�M.�>a�ր�-A�:8B�uha�\�8v�IE�'뚡���7�n���x��B�i���{CK���Ǟ�`��Q�	�	����kg\�v�5>�\Cp��\G�N�_���^���{�'�0v���`%̉�s,d���^� r,�䡃�H>RG��3�@L�ؖ:�4ӊ:ݬ��Ƴ�Z籗)X�HÈ�G�JH���!��+��Ν~$��!W�D�	V��B냅�Ӻ���jx:9<��N�~�N�e��ֻ���k�jZJ,9���P��H�$I��B�`�t}��w"`�j�5�C�I�@�U�Ip7��'&��U�]VnQ�>�If�����/xa��G���sY�R�/�
w�/�\��'��]���7r��J���$I��&~�,�c�m���GҴٷ�ʄw�]ղF'�^��=�Et&����y9M���c��(בW;=��ߢ���~���?6/�wu�U>;�9Y�x���|������'y�!1���"l��4�z܉�1NxL�\2��N5�p����,��Ѳ����]�	[N6(ؖhJ�I9!����|V'pը��Xh�E �H��6�dH�Y99v&�h]��6/=#�*��q\��͕c�ܐ������A�+�����4r�^�TB�-1Va���b(s�]�⠧�R�����(�!Gt�J�v,��*�4N'�n�è�͛�u}�����;�o��uF5�{�s�Qí���j�Fj��O�<�y������>|�<�y������>|�<�y���ϗ��PK   ���X�8lѷ  �-            ��    cirkitFile.jsonPK   ���X��2i  �t  /           ���  images/0d24f7ca-0a17-4a90-9ee7-368ce6dafe9a.pngPK   ���XB.7# � /           ��c�  images/1d5cef6f-7e1d-4016-8cd4-58d2b051ad75.pngPK   ���X����7  �  /           ��ӑ images/2b66d102-ef9e-4dde-8ee7-817842500f7b.pngPK   ���X#X;Y�  �  /           ��W� images/2d4ebd0a-2d28-4b22-8d08-8a7e71760a75.pngPK   ���Xt�ʰ
 � /           ���� images/3243dbfc-afd9-4800-9031-ef944cd75f6d.pngPK   ���X	�O�!N  �U  /           ���� images/32c80dc2-b650-467e-aae3-2893aaf2291b.pngPK   ���Xp�֣m	  (  /           ��M images/37476977-ab57-4ec9-9e81-825006455165.pngPK   ���Xf1:Ϫ�  ��  /           ��% images/385d3502-8778-4b9c-b5b1-c060638a35dd.pngPK   ���X~�`
C�  ��  /           ���� images/4249a833-ad2b-4779-932d-e559dc915ce0.pngPK   ���X��(�O  <X  /           ���� images/4b052587-c364-4d0f-a047-e449c1428d33.pngPK   ���X@��)  /           ���; images/53de0982-6112-45ce-8e57-c75f3734d94a.pngPK   ���Xwt]i�3  �7  /           ��0R
 images/612d2f36-6902-467f-9552-2a5db1e13335.pngPK   ���X�չ�k�  9�  /           ��(�
 images/76cbd0e9-fa13-4be2-a677-68c315f128b4.pngPK   ���Xd��  �   /           ���/ images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK   ���Xb��O  �W  /           ���O images/92294c6c-e025-4a92-b2dc-6de1496811f5.pngPK   ���X�^>1�5  6:  /           ��� images/9756906e-dfd1-435b-853c-fa5dc8217a1c.pngPK   ���X�&�}[  y`  /           ��D� images/982accd3-ee7b-437c-8e9e-7ebd1fcbf7fd.pngPK   ���X},��j3  �7  /           ��2 images/98e5030c-de80-4894-a887-e6b61185dba6.pngPK   ���Xǐ]zd� K� /           ���e images/99ae2b82-1d43-4592-a023-63b23200c4a8.pngPK   ���X��̋<I  }N  /           ��v� images/9a5024af-9389-4391-bb94-e3c02dff2ccb.pngPK   ���X	��#u } /           ���6 images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK   ���X*�x}�/ �S /           ��o� images/abeae39b-2976-4cf9-8094-7a1fdb96bbc2.pngPK   ���X�A�>�|  �  /           ��z� images/b5136140-2313-458d-a25d-eb2cb312f8ba.pngPK   ���XL�I�� 2� /           ���Y images/ecade926-82ba-453c-8c81-d3caca9f3c08.pngPK   ���X���
  a_             ���- jsons/user_defined.jsonPK      :	  �8   